��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��l�����f�J�éy7�=7?�w�e���˦��X��(|�EN��:D�*��{-� {���hEې�_�p�P�Fॹ(����ұq���[�A�

��я��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����y�GS�N>�(�3ҷo	�<Y�Hw6j���b���(>Vc���p��/u���}4h�~{���y=4��d���e$X5�rY�֕��g�7/�J��[�|>@��~w:^VUM���H����Kor;��Y^4��%迄��Ns`�_P�}0l<BA`�>�ăbL/tc� f�����r��<Z-M���-��^/�ŷZO�a�xI�a�"�I�"�`�� �P7l:� �Bz��v1��`�Gb��ϜVD����Jq�SHOY&0�/$�!�5uw"l���i)>z5!;~n�g7��Â��v̋Ѽ���(yuD1G&_�I*�~ԭ�hċuhj+n`\�wy쟴(���(#�3�i+6l���_Ο_��*��ט�����=��t��hH��"'��iL�ߞ)ܫ���+����Ѭ�u"��K�Ry��g�8¶�!�f%MD�<��	�b~i8z��8���cq8տ��%�-:P��~����+i��ij��W[��'�.������J��Z4��+�l/P��Åw�����Rv7:3�����j���2���2�]c�����5��L�aQ�mZ��Ĕh��>�i:�F<hh���&v�
��S��*��hjw��F����D�OYp���G���+�����!h����Ӱ�Qe?��93��ĳ ���2$mvY�'K7Ki9�����=�*���w��"R����|\�&��/rL�'c�R,��]at�ϰS(�N/r��e�d���'s�ݩ���^~�l��D:�}j)�"����~L�K���W�eC�n��֗�{ƥ(c����wm�ۅ���V�~��}��������TWc4��1sb��8��L5?���g�Y���c ����l)�D��?T!V���W-�R���ov��)X�Aha��-Q�����D���c�jPd��^q����E�/	N!\��w�1I��P��\��������(��'s평�˥2B��-	�@3p��"�-������8L?�hi����^7�
k��.fe>��1��G-$��#�)��2/^��L�?�2�3�ʩ�b�;ԛ���%h�g�ͱ�pS��#�����o�D���4�S6=�_y��+!x1�)a`3��!�4d�'<���ݕм\jҜ�|q��%'$rǿ��9E��Ѥ��B�^UI��!�(���)ZI�.P5����zuf;��*Ե�у�̜��Ԡm�z���h��/.��&@t����f_E��ξ����6O���D�!���yO-����pN
6b�fT*����%L>�m��n��	b�{���*^����H��Co�47-�*#�߷ٝ$��j�����a��U����.��Ѻ�u�P�(D�O����Z�2˺g)%�c�Z�⃌�&�S��≟W��H� 1�BCG����y&�3&�!��t�f�4�.e'T�L�|<�b�QWJ�����Iϋh��n5m>�Ӽ�ݙu.S�֠�����+����V��2?�e�~ۊ�uM��yߐ�Kڅ,�i^"�.�,��N�q���� Ila�<�X8��9�S�LEZ�^G.���w��O�OqRz?Q�Ң������$���oe&�zGQ�{���<�$��ɑQR�tࢗ*�JW�^B�xѥ�*������ftg(�$��'����AU��T����;U������k^N�ŧ� L��WHxK+�W� �W�D���E���z{��K�'�_Z��"Y-Gl���a�!)�� �1W�,�L�͖Ǟt�܅(�����ԡZ�t2�K�Ⱥ��"���u���y<"��ѢǠ���l���>;�l������H�����`]
��1��E~Q�_���'�zΩBT�Ҋr>�Þ����X��{�$������]0W!������j:l�8�4ǽ�ʆ�F�<)�½|��g�F�_*�#=�AR��S���j{$� �,�}�,�?����T�e�-�N(���y)��2�>$6DJ�.�-�/i��F݊0�$��(�d�2�bq,X�=:r^����qU|Ū]�_D]�������6)�>����Cdɝ�ʴ�����lj�P\�F�����"��X����h�S����Q��z@��3a�9���vr�,��� C;.�x���2G/��W �lS֊x��<���$��:"N�G*jt�ö��1�L$��r̀V:%���1V���q�*gT�C��e1\��'F�".��m$-���g�KB�q��x���i[^ӧ��V��-��	K�ˍ���(ڿ��3)9o��{7@�~�TR��Q�oG�R�:ҋ`�u�����V�t�)��]i�k���R9ڜ��'�C`��y����U�W��<�%	;_Z�ǪQX���gM:���EBt_�-��BO�)���mx���e,;v�UBOc�c[��Aʾ��2J���~�mڷ���.��bh����9
�Zjls\�#/��t�8i�N�r�\����{<=çjJW��%E'�������(�r���U�*�~���1�૰fdf*�1��Z=����l�y�����+� ��������R������9��o4�v,�� ����瞬p�Zѯǽ[m/�h�U�s���B7$��0,��ګ^P�I�b[z:ęI�*y[<[; %>puC�0��}]��o�����D�a��U��(�]��"�o��BQ]ed(�w�o�����k	G8�<���Ey'^F���Jٺ�	��p��>15*��4QPY�X��XMoMAK����0�@� '�9�C�v1�՝�j
����EKO��3����%n�`w�O���ȫFtxj�|YB�M�.L��[�����o*�9������'|��4�4ԟZ��ځ�U'��1���ԓ�n����u6
@�$m�97���o$�l`?U�� �aի�nZ��B�-1��@A0(��1B)�/�F�Vk���Γ�
�����S�`	"!�EL�&6[���N�:���r�31fz��9-��"�h��+�s�KgˤNX����������j�?���c�q=���sb!��2�m�ǜU�|^��x'/z.s6\�_�u�I>�UZJ��	'IT��,m�A��l�����ȏ�r�yrY�@���rlݿ�CT�M��!Wd�{�x���f{�����e�h3��T��l{f41S����p�߀f����Bg���q��_�6���O��֋��S��|b�hzq�M�s6;�P�q�<f�s�Ų|��Ҟf(\�������,���*�I_��G�X���B����Y�.���� ��sA��[v]��{Q�B)�|����`I�]�`Xv^%~���p1H��^�#���G�WZi{�����D��~��~�V���![���A��b��J^,곶�F<�#}>�hAf���{��T�p�3	 -����*^�g]�ܸ��O�Q��#:ײ����a�7�5�uP��UE��LM?��8Uf�=�p���a�X�EFO!!�Wf���6�D����_i�?�͠W:�3Nk�6�y=jMy��1�?�/̉�iw�����#An�����On�6dzx���GR���|�'�Z��
��sm��~�=���#�(��k��@��{��m�ѝ�Aǿ.!�F�U�6p3�x{{�K�]��k5%�O<�6J���sa�Y�
,iMjj��p��eW�I
��S)}w��yh��7k����Q�cxVQ�0��R��5"�}]`��
��C�!{�l =jd����mE��Z��ӯ(����+ӧ ��hLP$�膕a� Z��UK8� ��������IeR!\��&�71�z˾B�����:|&r�+ZE�u���%�I��yjI�x��-MC#����������ҠJw��f�
ф�?����
�s�4�9�ｃ9�U��A�2ZT�c�wzW�b���.�����@�HZ��4�D� ��x�-��A^��o	�`�i#�`����C�<;�����"9�7���䨴�f*��m���H�vtq�"�^T��)��!�� ^)�C@���2ps�"#������{�R���6��р^��eJȬg���hz�������<�T.��$0��������d���)���(}�"p�7A[e�7�V�$�3M`�h_�B~�1��n�@F�̱�ǈ-ڦꪞr�F@�6�ga{����0h�'��	L��ٳc�,��)�܄ޗ?ޔ�޿J�@w���_�h�B��$��}�.��6xq�h��*͵R���,�� ���1Td�Rf��C V\��1N8�8IO�āWSz�m�7+�&�b��h���k��?�O(��G�>������9U�=t.��_X���T�f�T2;H"�������!4��a��<����0V�9�eM|�ۆ��E6l^{c���F��8c�27��O/ :tɵs7�����	�R�U�����KuR�+��SX5AD|6~�=A�R�h���$��d0F.�=�Q�%��B�^P�A=`��c]i�$4�U����@�Qh���%�}�Ǚ/-���`�I)!r*9jG�������a��[���;p ��)�l$i&):�u:@����\�d!�;V'56.��lrd����'��M���/\�7�z8�~_�;fiW�<�nS������8 �jWB`Ն���Y��kȚ%z����R�͑;����z`�~ʉ*����#9�Ž{��@��Hɦ�t�B�I1*���(�P)�|�)��M0�<.���U�'�@}��[(YwX�\�����S\(��w27=���
oHK�죡a�L�Q<�3Jd�"���0�e�y`7g%Q}�
��ԫ2�,y��L���L�}���{����(\9{]$�{ S�]�Y@�d���Gy�F���%JO�^���nڭ��j{,F�?��Q�&A��bN<ݬ4$��(��ǁ��E�K���O?3wSq;��א��O�2��T�l�:P���}�8M���D����=�J,�
zAr7<���+M4c�?�ej�
�_B�ß��dY䎭#�hw[{�w(YJf�,
�!	k=#3C�&��7���^�^T���N�)��ى���䌵k��?����W��V�锪[�VH�4��a�ȟ�����s7�o�;E$�M'�ADc�A{�v�w(���|�&�Y�A4C���Mh�����CG��o��l9�0:*at��N��5��fT�Q4d���*��3>=�ŏ�ǭÞ�.�U`����a��=�U�0���od�l)me�+ڶ�<��b���WF�m�6�:���Mc&�����W�2�2>�O�t�տ�g�a���1���:���Tk!�|�eQ�8!{X�D�t�S[q�N���A�ȵ��dQ��|�<Ӆ	}�>�h�� ����|Tj+�����
;�'��>��7�wD<�P�'�R!�La�y�w��t�vXc�����m��go��5=�����%������	��g����[�J����e`����ۇ��͖�G�]�>ck�yn8����&A���=�c��\�`�R���x�DZ��
?@�ż���9ݹ��kÜ[��c�x+����ϡ�~��B� ��2��o�	�Yu�S��Ghl���p=mbW��w�u�[ j+�\�pU���|��H��9�4�'�Ix��<�e�U|� ��˱W:�hFᨙSKE;y�D"��c��{&�+�d|^��]P�؅�Z��`�Ey:#ܿW�~dN���Ya@���+(�p٘��V�Y����>@�=�^�W΄�N@Q��|[Q�`�8,��nՆ���b� �A���g�e���*Y�+��Wj�����#j|�z�%T�9J)��#A����ĸa`Dc�w\(�YQ�1@�Y�1�9�JY���sy,
�O�S�/�n�0�0ՙ�V�p�R�D�m3^�y5F���rvR������Uñ���]��[�R ��:#�s��rx#���̨"~��c��iq]�٥?�kn.6���D�+w�ʏ@AdÉ�HI�]���cY��j��v��1e�eo�� �4��\�+�g�NLv��@Uc����G#>����{J�(c���)L=�c>RK~�꠿Ne?�~����͉�#�~h���ߙ#\p�r;j�2U�Q�Rs����n�-|������Nj��z}}�f����o�?��6���,��U&�?���|��NEֱs��	A#j-�О5���ο�NQ3�H�05�fX���;�;� ���]d5��u�Q�lr��
��R�qq�;?��s�"�gS�%q���Gn�={8�-�\��ٖ
녒d�ơ3�o�c��/���i��޾O]����F�C?L��k����p�z�ly.��ŏ-1�U���K�*J�.���Pə`��+��{��w�w�{i�Oe)!3�D"~F�;��N4��֡�EJ{����V���I����7cZ���ULf�*|�]�s
[�ܾ�5���rň8�F8" }T�Q2�2LF��ǟ�
[z䪌-mg��{ ���k�\��E�G0c�0,+�r��t�ʋ�+��+����ꏺ&�}�Zj��UɎ�������<w/u,yd?~�F���\��f��F�Y�D�T�H_�U'�J�{X��`N���_#�-����Js��2sε�f@Έ Ո�����v;Y���f~?��~D���O�,8MLN�*�[�h�(��j`v�糣�u��y@��v����U�|�Z���<�o׎PtC���V�Uȕa�(*E��d�z����=����,�	�z�}����\�q��/�3���g�m�60�o�k����h�fsH
w�ےO�'#L�B�-a���^�l��#�Q��X�>�e"}�:��Iг�+�Q�����<G��v{�L�委��~�/+/�??Ƿ��5��N#�\���N�DP�^�=�m�q{����~yd��V[������G"��3��{�ᠩ�EU+F��2�7-��c#��l@8���uaӌ8U2k��9�<��w�0@6b/��@Q�y:��������;v����d�NİR�����@Tݢm8��_�~W���D�����bw%}��\e[���0����rM���xNkL��9�P��=����I��vf^��,Y�t���+r&(� aF ���oM��i���2�6�h�h#IsW���ec�y�U�l&n�ɮך@�&�J3:*	���₆�l���6��)0��_L���eJ�)�� ��tՄF`Cx�u��T�^3d)15yY�Y�#�$���!�h�VM�G8��%��Fѣid�e�����J�}l"��9/��ȃ��0`T�F��c�Fgu���H����&�"h���s��ۅ�N�l�Ts�2*��4m�fE�s�Y�7O,�z\ɬ�m�}fm�O��Ѩ{�O�.t�eQA\�-�1����2����T3���OE[6P_��"�[���,軙\2��vi���~Ȝ�Y�?kh�+W P "�����=y����=9N�@+�� ��+�\A��7ыM_���+�1Vp��]�$'p\��R�f�����l�������(��\Ɂτ�͡ң���Ͼݕ��c8-���O"H�=m���O��ݚ,`"�%;T9�躣�?�U��i�RF~���9���^�[2<B(�Mf̡u���.�<$�q��N�;ɠ$2b+bJ:��9a�'o�$0"빈��Mi�������h�����Qy-l�H��6r�0��6i�O��R4�/,��]tX��V߲�0�S��.t�J�6��X>޸����]�y���d�f��F=��E�,��~��z?7��0�l����A��T�.�L��-��.�?g� bJ�?��I�	(�y�y����ٸ��\)��K�z��O���A���x|���:��Z��7_�Pe΁hՏ�8��)�/@F����K�˾����K��86�7�7[5��c����~�@FY}�m�������ss�.'�[�|������M@�Z7��ŕ��{�Y"m���5�h�؏�8��L�\�K�j�AC�u��#��g�h>O�䡯S-`���_���q�އ渎D0w���x��(�l���~�}�L�-N��wE��<{m0GS��=>����^3ef�_�4/^�cȸQG2��A����)~�ͳ0΍�_������-f<6�Y?o�^{'���r��x��Jx�fTRN51���m�����H�NS�U!���B�{
ܬ�On}2�U1�YJ����y�"�<���ЄM�'�C�Z �A�䧑L�صF��L�BIS|���v�����,x�����d� LRzA��[:կs���N|�����p��>��_�p0J�T�\1$��>w�}L�!Ixډ�d��c�!֯i5F,��? ܵ�,I3L��L���O;����e�?��	��%�nf�����[NJ2 F��oo�a���c�i��׎<seJ��v�O:X�D���ӹcn�x��dͪ(	,��1M���rT���Cگ��`�X�[EJ1�]mO�0
�g
�0HB��5���0����{_�ӡb<�h��f�צ�aq���\�ݤ"X�|�7hg��1W}�K%���}���2���[D��+���j|>Z��*�w�<
9�f�)��y�j�!����~O_��3WWd!���^z	H�k3T1$i�K���E�ז�2Q��Z����rѹ�9`�M$�6��w���7�.b�F��ɝ��S/Ya�v��H�m�EH���5�Ua����K��e�W�:�Y�ff8�G�s#G���̹H峮�,�?
�I����5�"C�dg'J1U_�����d.�9ݤ��{�{��O�Th��k~b�&���f3���v�P���l#i�Ӫ�ai�������<:�Cr�^������s�����r5&�)��4Q~��'��}@��YW��ө2|3�6�)��Y���ю��027���٣gE�`��i��M۰k^���6GQ�9 Ʀ��m8����bb��p�EiLm���n,r>Z��1���g��Rٕ���uhu���}�ɥ�� ��%
KB��trO���5:w%xV:�GK���������W��4g��#N7|V:N�����B��r�Wlc�|09UU���e���<^w"�;�E���ש�Ee˳*�?�䳦<�*�.�Z���#Vֲ-,I?�h�N��.o]�m�ElG=���e��m9����p������sؑ�'(0��TZnX|�\���I�N���:��۫l@X�g]�C�a�|sǺ=M43!W%��xop������-}�$s'�!�q[JXyA�����[�]TCt|��DcNm�	���y��޿������%i�ĉ�Z���Z���!`ʊA���&A@�K9*6z��"��w(��H^��^@�_ ᨆ�bw ���8h��������h
.���jG��:��_~�*�����/���?�	$�I�`�g��z9[�Y�����q8r����k�	Q})�M3:�g��L��4��%l�a� u��ܮ9z��v�PY.�"׶[��
�6~��o�h���J,E�g�D��ԕ����X�C�p�Bj1��� ����#��ORb��a�[{.�U�ӊZ1ڸ,
)e�Õ��KM�I\���*fq��'�V,�5k�Kr�wZ�9�F$��E{.6�zlG��$�_X���n�7�@D�s�V��a���%Ni'O��G�Mi����%�cF�d��iB�v��r����d����[�D���w���WwgD���Gw������Ĭ��K<���'���4�?�u)-x%�#�g:2�|�!���r�/�)~!2�},VW�2Hi��X\�S��w{�ш��t���c�?]���I��w�cG�g>{�bW���-�.Z83���twף��Jg&�S�35�ғ	����<Z?7X����R>|_ʀoOxC�d�R��y(@50���h��IbI��g�Y��Z[�mЬ�-�P䗰����q)���ݛ�d��ߵݚ�� m��O�<m7���f�v7Uh�Tl`�0�1QS���F|�����)8�(�z�j$��g�K�F��l �Vy9S�[.U1]��S��x���"���:KRh@9C7�j�L>��O�w������U��T�ϭT�������m��G�˰�g�'Y� '�ﷀ?Wk���}���ȰQ���Z����P�t��
ׄu�)�;��*[��tw7�&z��-o?J�N�t�[�X9����fx!���z����o��ІB�V��|\�=KJb� &�D>�)˄���/gi2s�>�f��NT���$��E�0�ƪ��/�>�0g��Y��P��`�(,��;�{0�K������)�Qq|i�"օV$̿�p҆����0Mf�r�r�̨5,�ڳV����^��*~�:/�S^H9@��΃��p�+�V���c��8u�w��5~@�n�-f�%���zP�(qD����z��`���34+���ϛ1Rڪ�ү�iN���6,�V��u*�Gh4�|t�2p�P2"ӄ�c�ɷ��;��|�EC@/r�ӧR/�3���^�7-��r߬	�f�we'�Z��L��T�Е͕x�t�-r��뙺��Ym
S��j T}+�h�5��.��8��B���0��J�&��S���8{�o�o�L�P�!g��_) 9�E|�_`��w���Е^�%���h/��Lh=hTh�$r��HV=������2��"�r�i/�)�PL�%��4�!z�z}��hnp�|Ӛ>7T���G#��?	�%@�x@ �Cr���s���m_�At���Ikr4w�N}kQ K�H�@;�&��%B\. H�(��yl\BA�ӻnbgP/�w��f��)��������d�H����[G)�M��֘kM�1���l1k�J�&ê���\-�����7�8�Ud���j4�_��ǃ���ZT��PSCҺ��N�%�Zv�j+�=��:b4��_���>�b��M}i3m����B
٣����i��;���ca��k7f�i_�4OA�E�6�$�(�j�K-�]�,f���5��7����i�7�)�������C�d�F�5#I��˿�	"�+m����Ԝ��o�Gl�뜽��Pp�#�|iJ�{_���yn<�er���H��h�g���h+6p��8R�+����H5h
�cS>hm��Wnٟ� Hw��\�xU�-����!զ����Md�ej�,6T9�����\:�7hr!#U�c���3!�}�8��<rk��T5�#�.r�dU�PZ->��J�g��?�?�ߋ��(ܟR�8�M��=�R�f��v�!Z����*�u<�� 6�3Zt�]�/9�g�|VoE���&�Bߔp�d�o!�I �p�2S��J�NZ�!���;Mvs�>AD�,z��#�(��}�'���,5Vj��~[?-['�j^�Ё,�����ȈH��	ҩ����;��=o��t��Ω���>�u6~4h7���	�������8xE�I�[�>�0�����QG���{�-����6��F�!�L���ݞ�{���&Zup��i����^�lW"��O+���ﳾ�l�D�_����IŲ�]`<9X��J����*�$�#�� �0-��蜠~�#�U���<��F�5R��1�B�o�w��N?��Qz|��fG�����;��?�sD����@Y'9�(H� 3g�e9�1��Z����
U�ك)�1�ݭb%q����k�k�r�-���v��'o��ZJ~�� �6������E�[_;�"�i��>s���ǥ ��}��>Py09/�
�؆�ew��%8[5"k;���S�d�-�(?�ei�ܚ=L��P}�7x���I�AZ���ln$���g̿k'���3�'�\ j�*�/-C������_���R�A�{�/tq���,D�$�%��vlr�c&<����(���d������t��1���|Kv/�� # ��7Z(� ��#1���@(�&��kx����'d�jV��8<�G#�I_�����<N`�LX/�LK�8�����v���7�W��C�so�<ׇ���fV�����s8�b��v���+��킜;'e̭V5��#�α��ķs�:5}a�L�����W�xp�<�ۼ[3��ҁ�/Ł}"�л(i��7q5w�bJ���#`����C��c���6@7���]$��a)f'�B��Cv`�j�a�EH�P!���Y�ks��51)��q��X�/`�M��x|�x�ۛ�A��h
��v��lbF��b���P��+�O~����T�zpt�bm!��dt�G�Q/�OJ���$�O��VWwM�Cd18:�����)��y����5L�a��(lRF�5���a����a����}D���č�����`�X�����eJ~���̬{�\���D��WLh��.�OuӥjL�����Π�!�_f��$	hx�ڋY���l�?@���c{��7[R!	���p+Eت�N�ncԣ���<�Y��Χ0 �3o����vQ��"˜1��;�Ʉ�)"��w�9�dy��E!�]�/�C��Tz����yЪu�H�j�K~?�ԫv&<�6��+N+p@��\� ^���f���;�%iT�M�TuA��r~�چ�7�
+�;U\�$��15�����fd�Xw�Åb���l�9����(��N�0���݋ߞ�2	Q2؍�t��e���d��[�'q�����KԠ�!��v�]� �)�~�U�^�,l^u�Sq�	�aE������W�z�wh��f�%���o"]OC5
Z��w�J߾�&+��Շ��v�>E���H�e�bb[�GD�%�uV�"#�������X���2�{eE<�(\�V �UP�QRF�&��V��ôc�jB������}q�'�Δ�WXԫ��T�O���7�EE�.��.�������U�JB?W�~r'���!�k!�"�@�I���2ӯzV=r�9#�*�׿���������e�p��Ɍ�˺�{S:�G��s�*��C�J)b�*�<(˧ M(Pj/�[�L3�e��4�XL0��˄ò]�gEH/��B	�)���lE0L+H�D�2E"ħ���̻}::���S��ˣ~�:��r|pS��߼s�V��h<���*�����*�!2�-�I�o�q<�y^VO�m�8>�.;]e��!����U�,KV|����Gë~ t�np�Se.
����΀��4�ռ\���S�K���D-��S�pK�]� �)��A�3�F�>'�%�Q���0���G�N|�ɴ��m�٫2Ih�uwfp��,��=|m˺�]�::��m�8���y��{�J���|�_��T�A�J7���^�W�M�(�GMZ�ĭ��9�=d'���jR�k���2������z"�H�>C�w!��c���G�M� �#�(�oz�t�)���D�Cu��+�j��h��L��g�*��w*�������i�Q�����s�5K]����I[:�拭���������Ǉ'����j�x�{�3�3#���JG�)h�lEB@�d�I��������O��� ����(����.�H�'��M�p�R!h�"N7�锧�6�BSsR�+J�O�؝U�7��pc4c�hݛ��y��T�q��j�gl���\���xE�:RV�[7_�)�$�
���CJ�+Sװ��u,���ٹ+0�-����G݈�J&����J�
�W>ɛd����h�R���a"��,���ڢ�A;���U��h����$/�zO-0���ϒŒZ�A���4��[�_�\m6���ƹ"�t�~�L������=��Û��Rۧ�O��Q<��ھ��D�����(>k��\P7T�>|w0���(@�� �Fi��B2�0e��r:-�F�:Q�W���������6��xI�(��̙�"K���r��gg��#d�4)>L)���H0*~�<	��`�&gG��OS��K5��+��g�J%�;�H�`K� �{'�d3�R���~�p�S*���o*}U�%�y���	=�>� �B��$�����yW��p$��;�	]Z��H�\�_�O��T{��W���,���£J �k�0j�ս2���9#-&0O�K�{_*&Y�Y4h�B�}����c�4]&T�r�a��a4(�b҆��l;qzM����.�H���N*aD���QᎢ#�@d�ǂ$����'*=}���?�k��^d
�	p�8�jN�O��I**��-$�2���[`�\��ͷ�|�*ڎ�1ZYх�m��� {�@��H\Ca6���9NG��� ���nf=��ۏc]�%�di�}U�n��X.�)�d����)hX�f$ΥQ$����R>>Zx:�&D6�g`'��r���	*��)�)�ʖ�.������]R��u0��P5�&���_/�?�hk�#�����#8'\c������1�(14S�<����6�W��P.$H�� ��7گ�A��3��\[�����*[�E�L��-71X��R�ٷU"��X_0��ɺ�,����=�4B�D�s�%g{{L|8H������M��G9r��� �������<�Zty�|:E/)�M��+�Cd���8(�!�&�����(c�P�m_�Y��0h `9L�cu���#�	��=WÊ9�������U�o#�c{�̫_~ЃO�y�'������Xf�M�ӭ/�DÄ}���������f���U �SZ�;�)�dN��FIv�kUq��57c�������wV�ȫ��P�%���[/bF��xCz����rħ��t�g�m긼���	!QQ?�S&C�p'�?�V�,����(�'?iG�o��n��d�i�����zs�aݴB�W�<�?���Q�M�½�L�>l�sF���A���0<��(��0��qA�������ՙ*z"��?�	�!s���	�h
4 �<�F���(�am���z�>�ۍ���K��A�}0q����d˾�bN��'3v�f�R��')+dk����;��c��!�xۙ�M�� �{yxoѴh!��*qWp�h�~lxdW��� ��ѕ��UP���_���7[h�P|��O�t��0�G�l�V�i����¿�CkC�+`��- ��H.Ms3��h�Ih:)�'L�և-�W��4�w�Kݯ��{��#ķ��T�|L2*�Z�Oo4�n��|����Nt�D��A cXl��w�IR3./(�9�z��ý�\�k�Xw��C� RD�{c����J=�@��Ѽ��\#�#�1\�{ k*(�|FX`��K�bU�Z���S�O�12ƶG���lT�ū�o%~���t�v��� �9Z�;(����ՠCW�	Ed���{~]p��[����oo��04x	�9��H��J���hl���/
��X w��!X������JߋS<���pc��Ԉ��Z�ա�x���=�,\�Z�NO>=�S���ϩ�G�Z�#��|s�)G����U)1�i��Yw
u2.����Tq�E��[�9~���ٶ�m�`;�*�4����4�_�ϓ���71� ���~��C޹�&�Л���'֡�^�����F*/a�ҷA/��,*�6�pu��1��G�Q��f���q%�A����jOD���F/�/�,ߺK�:q~_S	�њJ4Ky���0c����.R5�O "&=B/9xOb�n��lo�Q��E;��,�l+ڎ�o,��sC�MH]�ϗ��6����l�� >s�_%�tg��j�_(�oɛx(d�7�_�o�}#K�Tк� ���yERD��s���9f��J]�+��>�k77�8���d�P�4/+v[�%�k�����a�\��G*NM|��4_n��N���-\"c ���,�3&�(�l\�&��0�4���ٓ���6a��W����ƅ��!j�kt��m睭�&f���j��F^�u�s��­�4L�HO�[��-H�p�d4������s�N�4\�(����=��#��LT����ƨ�5�+�[?Ґ��rGA��1Q���4�q>��sp�f������_������2Z��a���xautb��3k~�Zɑ�g�M�Y�o�[{C����77�!&�o��``#�4��� �aB0H��()l��z9	4��w>����0��5��z'-i�\��m�E}���{j ���wG��(US�]������52�!��N �k6�pX����5VG�ҫyE��P�VY�T곜�CK�/��[8d�{t}.nh��Ɵ�Z��9L�ZD�>��p�3�c;¶k1�������R)���z��������X�`/�����bͻ�W�s�	�0
I�ʌG�� ��K���[�r
�
����bA�aa��P���V+ͧ�fV��������D�����t�.5�ж"������Fwv�)޼��X��F��m������d�ɾ�Iv��:
���i��en���P�I���0����U����
d����;cn�K�5�ރ���:�|��oY�,Q�'�E]��E56������w��yw�9T�Ǘ���A�1��}6
�0WJ[#�6c�⨑nN��S<幖`�J�?�F����`5>�������_���6�7����ދ�|��un�ߴe��q��tɈ!(�z
#���IC�X���\�����������o��Y��򭘷���s�l���T��켥W�_f?I�*y�1��W�di�1�b];�t^I�w���7�N�1"�e�-��~F'Y̉����?�>퀟�[�׀NJ�w��=B��|+24ܕ�yw��Iy��2�s ��t�-zJ�հ��ʤ�'�=��o�.P���)B�ȅ���c��}彠�Ў������Z���T��	����@E�O�jC�>���vj����(}�(�m$�,i�y��C��b�����V8�P�Xr��L�N����������O�N;ca�,̱�oz@0Y�T���G��֪��z�L*�,(�@Y�̕R��A)ڪ��C`ű��%u��ץԍf��[\��I�h��kQ�EQ�245��֔�U�SqA���5f�N�&�W��fDF�٤5�����{Z��<�;<�$�
��~�0h��!��i������J�ʌl�ǻ�.���a��R4�}-+M�G���M;�Y$����_"Nl��^���Sz��{���*���祔޳x�|��V�1xb�V
P+貚-C��m���>�\Ԍ|MK����k�)=��_#9	uhj�\L��������[�z,6$���'�9�c��e[�*����� �kQPv�t!��t���g��������e�����?B������;�Rb5�>�u�+q8f���QGoqH�j��9�}0�F
=�=iy���N��PiIJܰ�Aei��"�NV~!�z��hJ޲�h=��B�q7%�*���{�~,�(�d��q_VVv$jҎtIK���♏�ݒ�߳׎��k��!��T(��&+�[Z_��^M�F�
2���T��I|���r�9vũD�LL\� Xa���bJ�!r ���NEuFO�8����Ls�r��E��6�����[��GG9�V�{���7..\��I�K�� �YQgO��u��C+qE�͜PF���ͫd\N}m]����wpLf�,B?2�uW=�)��?���%ցWST*��@`�xء��K�UG��?�^@�Ԉ�)1W�j91��j��0-H	���44����DL#M�lS'$��`�N�)B�M��;7���N�9׍9/ʂz�*�[ӌF�-�Xp|�D<�����v@���s��I�}��肋�Y�F[�|�����_�5���>{��~*s�΄�<�{cv⇿i6Ql&
*�;\tV0Qјs�#,-��К©ʈ�j����)#�hʺx�֍FkB�
f�4����"98�R�2~D}(=����|�;'C��U��:*���OH����i`�u�gP��J1A)���<�awp��߾�P��R��{,�oMiZW�s%�6��	;�O���/1�I	0�Z�>���.��[B��b�X��r$Nq@��	AO�to��
�b����$ޞ����m'YH��R�1�k>D�K0M������C�^�!�.�m�X]P��Q�v�ho�		���J%�d�CT�'�f�~Q-s�sk�2��>7�F]�u ���`��ؑdC��L����Nh�0!�L.�Gd77�r�c8·��B� �v�t������D#�8��� �v�ݖ���L[�,/xbؽ� }#����G.H���~�4hS�A�:C��;u/M"�ڀ|�5&T��̩1�0E49�;�{ZPѾ�q����-��=�[�#\��J_ �vʠU����ӫw �0�mS�֩��=D��W7�J\�F�+��)G�� �C�Z��?q1�v�Y'A9�p���t/���#'LZS.�K���1é�[4u�_KղG��7*���l�K�ȬR�h�x�Xid.kc�q�\������9�x�t,����.)EEJ�U腭�]/�t��zV�jG���ًv�y!z�P�Z>������D�ܑ��~r
���ĭ��:����UY��Uh��<^��V��Ip���3˭���$�tl�{irWP����s��<�9)��*W�����o�`�$��Y��v�4����,F�(oN�D3z�\�?%0���DeŁ��]�:ŝ��=9����#�����;ޣ?��/�ї���b�;�u`Sdls�4�YJ(�mW�l�لt�����$ƞ��/1=:6=�{>���D��Ձa�GZ�x^8�������*>���L�-�.�L����ٔ�\�.��L���%���a0��ϼ_U[\B~S���Z��v��d������6�J���UɋqrOA=��*�?������ot?�H��h�-��?v���5���
ʇ��b�B�)�������kλ~�� �J�n���5ް����D5:K���QO���NX\G=@Z��L{��,��-�i���ǟks>Ui���?����pى��t��ᮻ��� �q�F�҄!�V��)~r���C���;��o�`=��&��@W�9��lTM����w.��'����RW#�TMA3��5��ԉ���7Ò�$;���-�4��H�xj� �&W���<����RR0Z�����
X����������iG�A�o�w��2 ����[���Ϟ�P���xdCﰪ��N�P��aϱ��S�F�G�+��O:��ȝ��S9r��yk~�l��``�{����~F�`���rxK� �Q�8�$s
��JC7��s���g�Y�;�~�A`����AWxr7G_����'�NYklo=ς���q_�q��H��DN�@D�G��7�Y<���V��ǩ0�܋g�$�&C1�u�X*k9]3���5��;���70�f��B�n�l�H����ƒ�n�A���k�"'�ܛ����G@5�񆫓��˒0��#x�ԩ�M�!1�p���01N$���6���ɳ���y|U�����~$H8\YU6���̋o�JB~��bQ*��k�GLC�,jB	x�?䩱���Y~�i�ژȧ����'lrE����ԝ�U���f�����)��'�1��:��+ �z�Jo��g�h���EM�D9(]"������hs��iO-����m�DZ����,�Q�"�7%/�s2����y'��<6
�p?&�_���s���Zw��8q�μ~&Qu�<8e��K�!*�,�Q̷]#ڔ�qM��?kDBB�x�"��/�}�E�L�5�8��p��ړa2�%�."$5Sw򦖐���ͻ{��I3�Sz�.-ʑ�VW�Կ�9�o˷�p�m��Lʹ���9|�vxӖG����M���'�����K��w��p�X�β��ѣV^¾�T�I(uZ���
�g=Y@"�wP04
���$�Գ�_�ŷp�4o?�{�s
I��U���+_^��l�&y��q�\�B��J��ڷ�y�)�N��'��{���I�&�� ꮲ����A��w�	:�p��Sw�±!�ם�[������+b+__��$����w�K���2*.���� �y�M�fS��:g�3�j�[�p�C-��B���I/֥�f?�?���w(��H�6�={L+��p�w�:,c��?)	u=5�9qn��g�-/>g���\���.��e��YO\��#��ڍ��U�3��
l��[��1��F�����G�G_�+`�?)K3�we����	S/��p϶b�:<@��qE��:��@�.�����mE[����c���%��^r[b�fvy�FH1,^�T����0[d����?��I1����@z�~/��YRt��l�=�����b9�pRǾ(>c��@fՊ�s�T�	KI �4�6:�&��lj��¿���`�.#n⊶�k��m�c9Y�
8� O�u��]�s��w�Ք��!\�4� �qh��
�&�FQ9���?��[x� #��RF�5Ң��rJ��rI�\�s���s'⑋b#�#��L�r��q�L}Fu:�8��A��S��oq۷��b� a��1{�L��6� ,�Т-��?|❏��O���q],x�M
#ܕ�r�f�Ծ���n�@�T���k�fY	��;���`���P��_�'U8����f�����;�Q4c�g�a���@�-����I6�#����HÍ��z�WP���;��ɟ~p���<�.�ze����q>��1�\"N�=!�S�d�or�����M���Xr����W$�o���e�Ԝ-��JH���	��ı��3[������A�XJ`�U7��p�I_{L�J�?�;��k�"z&q���|	r�h��a���5�_ײ��]�d�H[U|2��E��9c�R9�F�W��K(QΝ�b�3��+_�qH�D��H�����qT	%͉;���5I�¹��3�ז��i��I����WT��g1��|m�6�Jj&r��:>Vh�b,u	˨�oyt��%��� ������&4�Cf9�!é�m�G�/�fG�!ީw��!��!( ��DO����h����|�t�a���<A۷B{�o�mf�e��M��5@$�j��`�)���+��,�����Ю(�Q������s���3��A��q�
���yO('�S:xQrZ�z�Yɒ��ay*P�/fq���6� ?NZ��KXW��Y����6,�/J9��m/������p\�o��� ����"�[6����Doe/���Y��aq�"�{0
�M6D�2���m����ʿC<Me���"�a�S��XL!�j��U$�����{��E^��j�R��ig",��w|�򑭔����I�u��W���"@i@ ��j=�f����@����T��0l�C�j���5{=����j�t�M���d?E�*��O�m����`1nO7��ʇ�~u��]�����GyEwEOr@�/�
mH��#j�с��SA:��O�K�==�w��M���I�qP���u�>�j֐F�KǎI@.���.+eD�.���Q��T�|U�;���e�=�iF�/&���'�d#DG��Z��k箑17PF�8���C��K��g9ч�����e�<�$��P/��>�A���*0�2���뚾�x��䟗���9;^�S>W�Q)�Mml�#���ܬލ��VY-1/{TB4>���^����T�&*�=�Y�c�����sOR�P���F�V��y�`�U��}�s�i3_�|̦lu�;[��g�6���rk8���w1��=U �A�A+��q��C�,���^j�?�a5u��(B��[��UW��pj`�h)(Y�ޢ5M�j��n2�ɑ
*��9#�p���0�� (�x9G�����Q�X�G7|2sN�=VU#���v��q��V�j��Fh�U+��?v>���Rx]m�&a׃Jۮ(p=����T����$dTpoj���}����U�o5/i�%XIqG?���{sv7�P�'�m����zn�^��d�K�I���5�/E�ƥ �g�l$P;]��8�	���Y=��j�>� M24r��%���ܖ�I�x$�i����^_�:�.�/iT&�z�����v�+��P̍��	��n�M���������j��<#��E喖͎F���
j��P@�yG��m�X� ��y'Rt�C���sC�K�4o���k)o1'������>���I�V ��!fL��M7�� �=�_Ί��L�<~������;���E��V�m��d�V�.Qd������3u�F�Yu��V�O��G�34aod��[eE;s#���]��5]d�ؗ9��r�ScǇO?c>|��g_�Cn������>���EF�dM��D�ZAQ�ݟ�:wvۡZ������j�������O��r?`��*| �^�<��:2ql^+ݓ�y�MO��v�"E�-&C
fL���~j��/N;8����G�y1F ��{��p�CR-�-�V�*�cZ|�����(h%/�M�-��G��H�qGf|�����t�U�HdJRy����/��>$
�S<���!�����ʺ�-h�&K��
�8O{r�V��á�I6�NYϞh�]8�Q2���2	������!�;	��o�	2�Y�����j��]�GG��q�hֱz( �k�۾	���r_����v���%�wual�{Q\�4�<�&
q��]����i�v��눦3�j4�)xj�d&�8޽L��I��S3�p�J�$AYv�v�4��bҒV�D���6����2�(_��ca���I;Պ��&��b��K�]�;@3���n���q�"�~C��hA�i�v�C���31T����<����P���������Q)l�拲E��!��C�z	�F�Mb�^?�QGi��Wi�� ������N��A���1��7.�D/�l왡�� rs�/�Ӥ�j��$��(�/_�Kf����5�*�9N\ x(�7���O�	��;�AP/$�`I��!�u=��5�TDݏ��EK4ρ�$�u�S-�nŽ��k��gZE�u��$1E�n�5u[-ow�`��X��10[{�ֵΐ]�=v�h������6o�Ciݑ��*L��h���<�h����8%��xCS�i;a)��}�Ϧ0E���W!�m��N��s��������F}�ml.=�f�.B9L\�m�m��h>U�H��ĥr�����u�1��ua�G4���;�'������G.Y��"��J`ݴ�z�P��	��?<�����.��1̵',�U���:�]?,h��y�9��ǚ��TE��ۚ0q����	/�Z�FB4B�J��V, �� �L�nR����.��������C�Q�յ \_�2_�����M�i0�ĭ�u������j�/A]���gd��y��:#[S*����lt)rMӴ+K-N�Q��ʅX��M�1��H-N�b����g] IF{@����[��5i �|ο��8%�v�����<8��|���Y�Y[���)�Ҹ�޵;w*l .S)��o<��&��������c._˶��p�Nۋ�^����H�L�����덽����	4�"�N[E����P:U�؄��2��'���7�Ѻ<=2����ͻ6�~	�Z���	�e씏��&?�YyQ���2�����.�%~k��ߓ2���o<��ϒ��	79%��	�^��Q|kȍ'h��>-�6I�����I��LS4'^��z�X�|P��K3ͣw�ݽa͚N���$+��]'�Pț�}��V*|�{��Y_���=1�#Э@.A�-87��!��ea"����j� ��[�_'3ŧek:j<�z 7�6Ua�hn�I-8jD�vߥ�ܟ!�Xү*�:��3���%�w^�y�ȹ�i x;C6����c����t�#�NĪw���:	�I,���yLf?Ǔ�s",V�D�c�J�5���ޙJ����tؠH�F�Y�g9Io^=��2M��6�$�|	����r=��Jۄ���,_�?�cb��K ��FA	��A8��p�>Ϸ?%��G_j�;+��8��z����+,��y;>�S���v2ܙ��תo�L�DG3�Z5��K�F�
" ����4�J�N�y#Ri��D��nk���N9����2��_�y�ؒQ/~�5�@W�rϱ��:�:����و	�Ơ/���,��z�a^A==������
�2=J%����Ϡ���_Ɵ�
޵�������Mu�Xʴ�Z�ŋB�̖W�2�_����Sp�K�x� #�	%�= ꒍j���F�n�.5}lh�_���}bYM��_��S��Q\���l΢㌧��{�;s��1���t�e�/x����oU�&K9V�UD����v|�#�|ݝ�p;�)���|�n���ԧ�1q�����H*i�Cl����!O��'#N��ͧMU��'�9Y&� ��rH��>p�-�5,/{�<GeR�ͭa�:��_vro�?�z�'����/�_o�c��VZ��r������b�C�-hI������GkQ�(�z���#�g*O�R�7?�{}����_a��8�E�?�b��k��T������ٝ�9\��F#�z��3��C�у�R1}_D�(o�\�r�u-A��u�W�`�N���mQ��PVB)���*ց^��2f�a�Q9��rC"���~ԏ|���5��m xE��n!/�u%��9w��OCxV���>�޻�p������|ֱ�YY�h�ge��M��-���À�텱RTO�5��<9%�� ���9�m��f��z���Re����<$Rh�B5D�GV]���7��kϨ>���ta��(o磝��
��A��\p���ӏ>[�X9���'��4r��ށƃ�0u��?��2[�[�a�:^Y���M���e��U��	Ȕ�UM1�9!���}u��g����a[�)a'�yR2��_[��d�x��|q]0�����_�ğ�U���i@ ��YFH	��v����9��t��<���Α�r&W���sq�[V#��]yf$�&U�����#����wS��X$���?�[XSF��Jך�����v��P��3����!���O�}u^�v�^��3�x�Z�T_PH
�	fUϢ)�/ ��TNH�w@ʋʸ`4CHǏ{�G4%�Z�;�JNVԄ�lGc	�zu��h���u���ϚY��6&�fi���<ye��/����wGm����@ <��,�ie� �<�j�j1�h�+�^��6����ň��W��7�6:d���?4��Ah
ʔ�t��W6�@QI`}!/O�]}�I�mJYp���R��w�\��P�Z���C�����V�)���T�V&�nX"�����_���+� >p�8,�Q\(���ų�cJ�5�@,�̍�TX&N/xUr��z"����|��FP���l��)�����L��pl����ʁ%M䫔��ݫ��f{��XDBU Q�TTW�D��ީ4�S�؜_�t���=y�cq���n��Y�gt��u����V�":_:c�%�߲����>"��,�����⨫~k�-��|�s����v���d��WZ������=�&鉧�{�Uz�+����Y ����,��A�A�Dz@|�(^��^ԅ|6�K�Fed]T׫��یx�[ɢ�*�s�ъA�L=�X/���3�4_
<�fx\u���2�t*�Z����^��rz�����3^W�GϤ�%�#�e��b�zG�&8�~׿�Ï�pO�>�K*|/��n�^���L�Fi���CL�!M�i�����O8�!��2�Z��[dpI^y�S��feDb@��Xk��$qgK���Cm��^�Zن�	���S�DZ�ձ�.]O���L���;tʠ`�L��tI��?�7�h ���\�KR_�3o���^���nz����#y��8.�3�C�y{�^?�yV�sܰ�S'���f�	�\ޤ	6���J��_�s)hbR�8���� ��iC�$������[_��TA�
��+{Ns���� 4�U� hͨ�*k��X�#�T��9��W�˿G~����}�:�-����_����BRF�c�L�*���)
[��fw�\7���� 9��h�B[�yˑA=��Z ߋ�� �G�#Cl��l�/;d���S�R�F�E�pj�puux�����g3��㹆e�$x�{�Tl�[S�sf�_��*�rR���L�7K�����a@Η��[�E��q�llN��h��gmD�B]�M����L�NQu�}W�6�^�4�2ߖ���H���M7 V9+�:%;�[�Max�/�p���v����aW��[���$Al��Yzetx�mY)Mm�@�f��!`A�k0�`��F6�@��7x�����j��k�B
_1��i�N�.��jȻ���hq�&��O0U��v4�j�N��?�`�H? R/�%���.y��L�2ǽ/@>d��e���g?t�.��|+�q#�Y �ю�x�c\b���q�4=��@���&�9Ͳ��8C#�.�R��ٕԎTTgr�UQ�B"�9����}5A5H�s�8V�ud��{)�LtDXI�:�)�� �����v�3�"�&Σ��)���SvBZ�:錇颅g��=�7������)P����3|i������zc�YR��)-��>`AO�')~�2=Q�+�!�N"�28\��5�C�0��"<�w^"j�XDB�&�����w��)a��W>���w#|��<���F~�j�^/��