��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��l�����f�J�éy7�=7?�w�e���˦��X��(|�EN��:D�*��{-� {���hEې�_�p�P�Fॹ(����ұq���[�A�

��я��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����y�GS�N>�y���iȨ���?<vl��S9ׯ��ˍ����ܜ�eg^�����|ǧ/XgߐB���Y�#��n�ig�|Z���X���9�
:�dg�"/
u"<~������:zY
�z]X��Ӑ�#.��#��ԅ����-n_��$���ܡMJ�l�����h8�͋��x^�k�ڔQ���Q)�p����jy�-�PTh�m�tS����>�f��P��d(+�U��,�����J�S�x���pױM�PeP`��&94�Fa�c�5�rT�n<\;h�msy���K̙N<���9G���K��xw�����!n!V�]e�; T�L�v��^vT�^�2O�W���hœV��1;p�pz���ز2�[ë��L:�]�lf��� �j"B M����c�~�B��.��mrr�4�R�њs
ϵ�*q���몕�Ҿ��ߜ��Q	�QCQ�D���y}�݆�n�pJHc���cJ�����Dn����hC�|	BW�p?Cs|�_Ԋg�9>�|4O�j�Ef�vY�&��H��6,�KJ�D��8$����_���k��H<X���א���A��j~��5/qQE�O�%�&�zV���t�BM���I_��ʙ�v��7�^,�|�%ͧ�X�.�XFA|�0L=.e$���� �3�X^W��4!55��պ>�?S�T���HQ�.�Q�xs�M&�/�i����B�j}�M�t�}����,�3:e��:Od.��hJ��ypj�_��H�жJG�0�L�L͜�k��T�/@jR�N&��GO�?�	��S.�j��h��1����	R����uL��"a�2�iQ���V<���.���G�*vU?������3Nn�غ�4�lh�%΍�� ���|��� 1�f+�T�%��Z��tI9[Y���%C�~>?J�1L5Zp�_���:����
��ʸ�2Ӡ�9�hF�gSfp�chX^�cA>k0I�7��aUU�f���&��gDY3����2,��^�n�	��o?]�.�7$�ћT�2~YM)�hV��"UɇV�~B�6�AK��[ꮜ��H҇_֏�I���3���xڇ�l���TD�ׁ���l*�t���L�Ȇ#�&;��`mD�˱�qy����~�6.;
�gԟ�u�4��7`UZ_�<��Η:򓰓v����ѡ%�L�X���5��ߝ7Q?����Ip2�2�/�u90w��t���Bh�EՀ�i0t���?&5+4_`��Ň{MF$�K�W�HȢ�'���9\�`�<��������Z���0���3n����bʇ�]<F}�O���k�/Х���f:u����^�U�k$�^$0�B�V6�/<�/�f�/Z�����=W�Œ���m�iJ����6ؓ�`ʮ��L�+��m��ő/p;>���ACHlm�L)"׬"�B+���"�h���;+{�8�cܕ´�R�2W���'�L�k4��V��
�N[�fӰ}Y#�i��\�{��3cʝOÁ~H��X�l�Ӭ�y��9e�v�(��Ӿ/��^ݡ��4q;H!�A�Ђ�q�A|s@q�N�!W� ^ ���:I���P��������uX`hT���H1F�,�|�b�!����<���O�>��jXMGs�0x��H�$Be�z�]�ߜ��J���sy��5�0q1]][&���Yf�Q�4ǉ�S���8m��$�£M���h�[���G�[s�H����˅�p���ո��{Go	e}B��n��Ĺ��,
iez�0�X{O2�n<0�v�\G����v��¨l��<יAY^�x�h
�'���!�J�_�����[g�^��a�A�D��U���	�.5�m�yK��6��Yxb?�k��]^>
��$Q>/�����B̀X�!�u"�sn���"!��,p��p�^�p�uœP��>S m�xw�����Q-��ɉd��ǯ�Z$��-�����{�?b|s�5J�dz���VT:<�Il�@�ó�.����s��QΝ����obt�|�Qe����@�8�H�?�B�T$���c�����8�mӉbH�Sm�8�")-�-��@�Z��H��5�j��Qr������xc�8��.�� ӏ���		*.i�PaN���e�C�'�˩p*��2�ئ,9\E�h�D�)��X�g�� �&؂�bR��3��I��~x�.|᧠L�#��a�4��Q�(��'U%Ĭʬ��S&��k]
�F��1[�b$/��j�Ǐ�ye�5��5��w�������Z�v>�#o�
g˵H��\��7l���k��|���EK�c�@�D@pY���,�M�I)�W/+@R�~�_��9V)gDw�Ѝ�K�>
����]���/�L~�)������ f)�RsZ ��5�@ P۸g�>���
����mcM���v?R|1�E��czx?�]��6@����/��n>~ch�����gӕ�sе�k�KƑ��\'�Q+�	Ĩ^������e��_���J,�5���X�5���u�LS <=v��[_�x��� v��B�e���'����3�̄���p�?����	�x��4�㵶[Q��u?6Lj<)�Ǭ0DqM�Hq��	G*��A����Z>�ՒrT]&C7�sכ'�餐�nP=�nW��v\�n��>q�9�*�`��j0��?9�ޒx�:*�ڄg�<�u�ʟބ�5���F}w���� �|�3��DڥQ�$M�gc��ysK�M��$E�EOA�� �{;�56ʂ}��
��yǌPc���|�g�*�t ����-_��8k*t�j��67����0�#xV�.]"�E��fi8t��w(*߻���U�͏M=�R��$͛�I!���+���z��?+G���jBږ�%KYj��'��u2?�=ՄW�m
r{��ۣn���\�I��Q}�ޫKe0ܠ�t�q�PV����˭>[�J�N�+�N��Z�ۀ6*F@�����!���q������/X6@N�I$��X��S�5,E�~��ј�k2"S������]Qe�Y�곡zD2�d&?�vZXh;����y���d���^p%Y�����kU�nP*�7�rլ *4��0p�7Z�v�����"�A����ҥ ef$���Mt_	�hf��6�b,X�lP�}ۻ���>:{SiO���;A�IL������9�g����;j��A�E�	���i*��/ޱPMNQ���8��Cp�*ׅ�N�s�L(lٟ)�>އ��.V��{-�ۀ�}��D�\�a+y)���I']�"*:h�}��V���׼ہ�3���-��t�F\b�y�5��gʸ�����������d����f���(�`v�wW���F;u%�1�B�0H��?ı㕏ι�����gM�H�J@���Yl�d��Ks4����oE�'�|W������&�-��nG��A���+D�K;}q(�ڭ���&��d:�q�q��GJ�W���Ղ#�<_��;��҇��Yy�_}kƣ�q�#o�c:/��+໰��F���|�YI�v�>�(*��(�Gj�g�%�q�/�����5���n̓h�����K�J�v�2b�zŠ��9�ȻPo;c�Eg8����=�0%��VҖ�r�ֲ�MT�=yŕ���53l������l��x��^$37x�Z�F���T2����1oU�]hřS��)��=K*�ڑ����`>%Q S�����^t+￻�"E�QϟE�W*+i�@���ti�P���5E��|�T��҆��;�Ħ�
�p�FXܙ��z�[�84�>���(��e�,"ɶ�������O��XuS�=KP4/�vྨ��u���a������]�@_e�$�a8�?�b��T��b��pY
��s����8d?o��<7���A�,����]�Jo�v5��0we�-�o�la��i����@)��Q��u{�񋷘 �K^��#��yK}|��4T�&�&��G�JE	��<����� ��A����<�2捍kW�a�3F���us�m%Y�^��Sh�����4?X��!���0��z,� �HzK�X{��{��g�$��n*P�����V��PGw��N��y�R�ҋ�Ϥg4�i���%��� �K�j�H��S`Y/L ^�B^���K��k���x�JXAox��$�E��w��2������������O����O����!�$z�!^/S���;�� ��dW�:0?t&`[%W]���vw������+�"�\�G����E��W��IU�vu7�nǁ� nl�ʨ�O:����q�)�H�����n͑)���61˵��!�/��9�w�͛����+F���h��kd��E*i2��y'������/`lU��Rvى�;x�7Y#?����7tG��}�A������d��ɹ��!V�)v�D{��K��Zjr��h�_~���05eS��M'�8��N2s� ��z����=ar�&N�4J�p+N;�@��m�h�]��"}��os5�_�����L9����TԺ>��%-���$���b�e�����v�ٚ��B�M'�p�Qgcߟ��&�%�e-�̌���,ۥ+v03�D�����,p��K%�~���@h;Eu�dk@�U�U�yT��q\i�Q�z�:��~��Y*��8�{k/3��,Tlh�S����Ⱥߋ�=�Z������8�����c�BAE��X�����rA�*U����Y��}�L(1���ig��m"�L&=s��3�xY�ktg$� '��wa���ӊqa�]�bH��˽�93���y���z�]a�.�0�~"�x⒆�S�	�t%?��0��3���]4Ϟ����	UJo��n
�K ��J�ˆ?��`��`N9�@��q�m�{��a��V�a3�^M?]T�0�k��)��oQ/a�P������d���"*�i�����E�$����&oC"g�|	�rB�Zl ���p��ak��ԗ�?�qx���#U�=O�@�fkʁaR58�%u��B�12,���q���^�1(T����_�"���Ag?<a�orV��X&�v{��I��E�:5��p2`e���S��Cq���31��4A��z���6ܟV���P�_��I3I��Vs�y5��|K���%�Gm��o�U�N�[P�e�>oxWo�Q:[Gw p��boE�{F�!�5dUc���2:����h�F�u��-�g&�?C�%,};�Pˇ�i��Z�T�n�Z�S�f�]4��Qq�5]�+-��!D���*�&*����1}�h.d�-Rʗ'�2ti��Ue�Z�U�5�;^���$�ch�/���rD��� ��Nܗ�;��4%#��W�۪sA��]n��|`5@��>��,�l������]���9��'��k�{D�c�(�v��t���b��Ǹ��*b����"�=�HFv;.�NZY�I�ߥ��|��9�m =�]�����O�Ü��79�:}E����4�Y��~x���""Z`i�{�������a�]���r3v��ިYt|S�j�*��p�L����\�8��m�� 5��;��n#�%r�%X��27��]Q�ң���'��$�*��y�( � S�J���-WL��L:$ab#}�z-M�ǳz+N>1'����������kH�EVT��Qq@k�9�!Sb�6��s�A�[�<t��?;4���]�a2&ν�q�.X���A����q��R��*I�/$�/��-�*�]`���Z�ab��L��i4i��J����[�Z������2G�ڑ=L�7\G���J�5���dv��w[ʆ�s����>��f��b�R'P4������^+�&`_~c�F����;��G�x85;�j
vө��}Լ��W�3U�r�k
�#O�cГ����y������8֫#SE���`�C��`*�����`�$��^-��� �5[	�B���h�PjF�_��y�/b��T��,������\|�#�AnM�D���`=#��u�b��Q�B�7o�^�+a�@;yas�	�K��=ȉ���N�m·��4��Z9=��7	��.A��
ʨߺ�ǭL3e�4� :�g�&'��Ȫ3ů/<4�H�1��۹��Z�A�����?�D�5<�O}oF!�A��k�
P�̤;�y�_��y�A�Ű�R�'uw�5��-���z�?V�"F�'+��A��#��>�9'�zw��.0a��LM��ӌ8����ݭd̷8�3�$�Bx?�C�TO-�]Kr��&�D�/&��R��wv���D�c��2r�A���j �%�+^�oA�;K5�9��8(FR���1�� �\d�/�9#�7*d��� ����!L�(�`�uF􍱸��iB ���kLgF�"Q���F<����[~��8QR�_�Qu��I�)W�k�E�q1*�B���j �g
��3+*�#�3�z��d2�pW֣5��8��=v��l����V RɋL�=�±��ӷ�Z4.�����d��׬@��dO�h�O8�mb��i=�ᗂ�A�P�Db�n�dh=[$�T�`&���u��u�6� .�Q�g�W^�hPH߁i� >��_�ҁ
@r�r��6d�C������	Q� 	'�X0z/���M��Hn��ֶ��Dd��ӕ7쐛8a�M$#�+��O*��x��"��'���E��M�2��$��o������a�8Dh5��4(E��,w,��{�U�8��0q�s�K0�i���"C6�~"f ��|��tpl�6��ל������7��ΐL$�7	?�H��]��L���r��Aˮ���0��]�^���-����V�^h 9�Xk,S8|��s�I��f�aX�L�3(�/�������2k��)w���;�'L��Z�i�<ڡ���f�O�0��*SOe�7@�!Ӌ��z�3o��7g2~�_P�X%hRt���P����>�����*xg������={f9�`�(5�@��~�8��	�۩Ն� 4��Lq���"O���$�\Λ9�BM՘5R&��s���R`�J���W�0�0V�_J���9E3�/�#�55p�aO����f#U�W��u���RP�񃌓�q��}.	����&|7hɏ�Wb���WN�K��$nKna��ۖZ�u�δ�P�,d��9!F��rN=��I/I)���WM�$a� T3��N�	�)�T�}	�lcG��{��D ,�{��p�h�z�˸���S�h"1:�X��[��s�N�o8�}��������$���Nl��Q��ѯ<����I���R"�u6�j0͇��-�?����7m�2z]+��/d�+[=�nRY\��B
�d��SI1����&����C�u���]D�����uĪ�5}�i�7:2���<��Plh?dx�m$�0P����e��B��������pJ+�������1�!�3��˟w6�gP�"8(,��:���R�$���W%��e#�c�Y�wBx@�P�]��:>VK^���=�ħ>�x�o���E��\,�DY�x͊�KQx8�5$/��#��/��q��1����Zh$;R��=iD��� #��i�HD��\��@�N����O���=�?�h+�x�Ԡ��TyMTϑZq>>jK�yr����2/��II|q�}L��Xy���'���8�#ǯİ1��7υ�0F2�
N�^�4�g�&ũ�,�cZf�Vv���&� ��~�ݵ�`���ڰj�>�@�P�`�K֡������@�pN|Aр�#be!*SK��]��)Ue[�J4��D7������|�V.�k.��:i�����.<K��N����n���6�W�]��>�e�Q�VdMD��h��{D���� �G�	��.F$)a���EU����Q3�sUu��}ޠ�D���i�I�{7�0)����W�J���hE&:K�i�֥[g���o�V�G��T�4�?�@1�i�i"�� ���'� ���G�٘�F�[�� ��R�C�̢��+���U�w���i��r�1�!J(^��� ��e�n�)��D��t�q�LS�U�}��4?w����r��R��ᔙ ��@�um;?�y�y�A;�'�A��Y�*�#�H�q�sq�ۙ�����r���Fߺ��
ۙo��uzr����ӿ(͚���+~@�,�<)< ��7�5�'�o�A�6�3�3��*;�jEb ���<1�(�Xɵ��v��*��{���z8�R���{��}��(�)	�P�ɹ�,0�;��-_���U�BAɫ	,,��KH��o�hg��w��;ԕq(X�����OtK(�raK��}��!T���,�SP(s�x�¡��V!��зs�JW �#�2�D+��u�.$~q�S1�{r���P>�?K�5�|���jS`��i{٭��@4cE�y�P)�'��T�;�]+�l:��z��Cu�1p�*��l-	>-Daw4��+�]<���]Mݽ3��E^�¬�k;i�+5�.5p#V`��!+F�lv���QG�Mc;@t�Q������������H��03!�Ϥ�A�g�������)���SE�qn-b�$��:������2%t����F�&S=���q/	t�.�����`D�y|�lN$݀akMۉ�,Dx<\�ЏB�Ꞑ��9^a�vh�����>�����}��t`D�����-v3�@�o����_{14:�Py�Rd��Co?�hO�ZKҾ|���!;y{"�*�P����?$�	��]eח�h�ra�
����^h�3�z���f�_������9�Ía]x�8MU�D�!Qs�2MJ)�AF��@M��UO��(>k�I������T��_�V>4n����n�;�4��#��@u1S]�0ݕ�[�Jb52��^���T�`B��п���jJC���H(�p��uZjS�fOoc+��D���c�..p���J?Ml2��?MͶ^έ ���� �p*�dLVk��w/��O�H�M{׮-I��m�����p�����&6�=��Zعު#��1�/�S��x� js��D�J��a�=q6*�a�̴��2߲�S�٨�^�<����*0�\�&�����ep(e=��g�~�0���HFL�b�h޿��������NnE]��9t�AtS`8�YŔ���Vt�>b5�է�����qKl�R�ޙt7{{2.�%��L_[t�X�xs���d�}g��xR��M@@'��ߧ��𭠐���Pu��OiN�<e����\��ˏGF�9*ZJ��`�"��< ����κۇ�QҞ�j2�� rKlܹK�5ʟ�񚺘�N�����|[(�D��V\w�Mzn{��7m� �^�'���'f����!��F�D�ϙ���as��s�)���#�&�W�����mi|�E=�mK��rWR�|ھ��K��P-��~9� 7�j���	�Y�׊�"�w9��\-}��=^���BG�X��/:X�޶�B���ux�5(SSwߴ��D!r�$k�I5%mn�8E�RA\c���d���ȋ<��U���U��H��E���K�;��T||��ʦ+��L'R��Ϩ\͍?��dK�K���}ɰ!������ڽK2�Q19��.�&�,���zjGi���}A�"��z�X�)x�R�X�W�Ź~���,d(���C�L��s��ae�FMP�^i��"�8�m5=?5?t�����~8-�aF�d�,�Z�byY����	���#y���aTZX�u/�uSڿ�ϩؿ�QT�>�!�^e2��RJ��T��