��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��l�����f�J�éy7�=7?�w�e���˦��X��(|�EN��:D�*��{-� {���hEې�_�p�P�Fॹ(����ұq���[�A�

��я��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����y�GS�N>�͆D�I���|NO�`]p\9Eʟ2�}��]�*��q��������`���@6k��{l�- N�c��&v�9.�\ɛOBI�{l�s>�)l��Z|��0��~���  kQ�d�{�]��9
r��A�X:)�
����>X;W5;����E_���A����"�7��z����-��\�_��"��C�>�X\�W���D��EW͖W��M�&�umrø�a�H��ap;~-�㋤��o��E�z B��n�Ŝ�vO��_��`�eծgE�}@7%c�z=�#]u��0�|����q1d�U��?b�N?>M�\}l�u�o�E��7�-E�{aR9����2�gC�8��Y3H�#_�$��Y��/r���(��}Nۊ�����<,���d����QŪ�4�,R��|��>�j�n����=��m�f���$/�@&�G����嬩��D�����g#W�ζM& �K,*K3��,�p�-c�B����8{p�C
�B����0tr���@��K���I�v�r�.�aW��Dep�I\ٹ!����{�1��S�iE���-�edC8z�X�L+�Uq#�d�V�z�D��[r�i���0��'�4���J'����qS�����Z���pj�hQsXrO��-���dS�bc־ï6*�yve��}M�x�,� ���|x������9,�ڛS bo�ЀX\���M\���v�Ob��Bq�c������w�ҟ��L���ͽRo����Ŏ k5V�~�s+��hin�-eA'ܰ5>���첫�H�{�#/�^j�ә�8y�;�D[!�k� ��{�!	�ɚH�·�]�w���$1]:�����5�����"���^J�A}�I��.�H(G��ʍ~�� ��.r{5�C�Ϭ��6���ʁ!�c���it�ȼ��y�n�{#�X�(q�ʍ�55��]y�kƣ�#)��O�  Us&P�2�u�iCU'p�?^��:ղ�c��$&N�}U߃Zw �Y�y�9��T;�;�k΂B>��q�h��B���ʒ�X��k�u�P>�*Y�R��,����c�C������$�q�����F�?�*��L��N)h�<���H�#z2�x�ԓ�T��߯;Q�>8��M�y6��V��Z����-�+�.l��Y�~
�9��KѰ�Bz�<x�Y:���3�۬�؃�Фs_��w�	d�\<6�ѯC�1�qCr��|�d�n�q�މ����2o�Ly,Pb�Y͸B��s��*���FЍ��x�v��t�z�W��x��tA�G�n_�w�0����:���f�L��,��C�P�%�{:_a|)6��-�r�`uj9��F���q�D��[`�0{�K��ޞp��v��Ox�ϹæwX�m_C�w�"1�/��-&�>��qB����l����q��yd3���n�����e}��YZ\��� W-%L��F��T	�g��dP�b@=� ��~��-[ r�W�I�h �61;�"��v���b�;¼~<Who�X���'0=����@��F�Զ��-��F-�U��׮ ����R���?#���;+���&cZ�Y\�m:�WJ�q?1x�0��=����+���u� P����Fk\c�i<�o1kE%BWT���
\/�-���ۣ�%C���U2P�.��8#i�s!G?:���C�*�e#�~��F8������57	�v�W �	rϘ����3 �����	�*A�S�m�.7�T��M��[-�g���kѮ�*�g�۾��"e
 2�n��I��ؐ�N�m�}�V��%0��lS�����	i0����
§Wm�e{����E���)79�J�\lD�� ����l>܇h��^o�!�WޠiÍ��KoA�9�^�EV��wԸ��}�v2Y.�4ĖF�~�U����� �;*��)��k��^���X�^#�����d�`�;��2�������������F�A���:�k4S��B������t�ŧx{H�*�vgB�ǁ�fgDG̬�/�^g��m���Z;����3�m�%��u�)���hb>ui6��
��M��5E��� �����-�l��͠؄֪��-;'O(�i56����O��γ�:���ӧ�2�5���u��xY[e�V��%@��>m=�s=w t�Wrd�!iT8�d�fq����g�H�4�;�zeŽF�7�@�%O���*h�R�'T�r�U�y�SO�l&n��G�f8��T��N����u�^v!ب~n������v}�\�M	W$2c)�^�����H���9�ݰ��gT�v��"���&�����6n�n�J�K�v3Y\-�Lqs��OM)iBl_Mf�u@�v��;���ؿ� ��p���A�rA�f�lV���j�G�*xV��N��{�E�l��@�aq҄P�+R�����M�5Y�c��żu���sWk��K�q6�$�Gy��/����31QV�}�GI����\>�T��rA4be�5Bb�����R�Iŋ(JZ�Z���I� �G�3�K|5@��d��E�G�ϵ��#�E�����!J� ������*u�ʚz!���"a��#�U�ul�O��C����B�2�V՘�B� '?JW�9�����(ꅦ!<Ƨ"!K�U�#�x:å��$�x�ri���Z�Jcu�+������N^�����j���^5��w���4\b��_�ly�'9�r�{z*��_���t� ����Ū%�j.Z����&瓵��w�Rh��G�]�Z���S�Kt�ּ��X�I�'��-2w����k|~cF��d���l�Tm&���`�LUR��7b���9S��Y������5H��;�vNf&�ױ�;��a�j(���Խ�!���08�4�5�_�Y՟b�]ʽ+ �^��b�m����mu�s�)T���8�gY��h�b�=����wn��}<9�z9� �y&z�A#��ě�l�>[ �X��x`�^p;1�͓V+�11�r��p8�i֎_�ex���KL��!�$����A|�����&ȗ���|�r�u����"���];o;�0r*��'VN�����j$�bc�bVP羑.��Z���F�؞������q�¬�Ny� QIȾx�Ro*<����7H��u�(�Ƣh8v���z4�PƥI쮝��� �z/��b�3䖅�`�N	Zc���S��☏��/g���=3�z���&��>m�����(5z������WĿGL����trۖ��5��[ڳ�]�����(D(_B�fǷ��L]M�R����hUe	�/	�Z&8�-���u$YwX#2���q�$�	�G؃���g��E��'�e��&YZ�p�m�l7]r��sy_���g�Vj���Y�nÝ��6_k!�|�%�q
�KUca��1�f��8i�\�:w��:T�� ����f�?��+��
�i#�a�ym��,�KV���id%�6�t l�t�����߽1S)�FKA��Oo��l�b/�'_rqHJ���k�!����)dͨ���H�\�#șHH
���� �(��F��*@�p���}O��� /ބW�ܷ��#~:�ee�u6��3����b%��Ͽ:��� ��볰"	�i�d���("a�j#�>�`]�/�C�_��W��&��;���A\�����#�]��ř�0��E3�ִ3~݊�X�^��v��k>�&ȥ����w�ږ���ںQw������	�^��֏��m�W�˥fý-{'��d�Fw<'�.s�2v���.�e�ɕ�S`o'3�U���ک���o����������ZM~JX��r��������8���⊹p"r�a�����`���t- �1�����s� ћ�=g% ����Ѓdc����AԂT��+/�=�d\�}��@��B�����qy����V�Cq$��w_���ds-�SiV�R8���B�ؒ�N��o~�Ϡ���xB���!~��x�R�핍Wyӈg�E�Ңa KbV'��c�?2Xܧ�������gS��?˗S�ԏ�B7!���C�-�`�9��^7EŃtF�)�%[�� �h�?s�x�#����?~l�e���΍�+<maџU��l���7�k�B����D��W��L�����������0E�X�sS���g���k���d��x�&U��}A������t�y0�}a�,�x�:��BZ��R�|[>�d6��S��-�	�9��ŧ�R���r,�E���}y�\0?u~E5��Y1�Sy��&O3��=1��9�=��uJ'<��K*FC������F6��I����;����m�"}�{]	�M�C�qJ��m&�N��}�@Zo�P�15$Y�<��p��.@;��ݢ�Yn���x��%7����"-q
2Uh�
'�_�6����7�ov��J�E5	�� ����� 8�L:.��y
�0��x������i?��M���ܵ~�fګg�Jv���.��r�����t�A�5�2�t��b�0OML���y_�,nFUX`��	ɺf���cie�ȍ%I��1f��^9!���5c�	��rI��<�@�]�`����k�>����j��؀����ʻ���'N�q��eO���+x�Zg�0}��Let�2Vb6F�0H���²�����Dsf"\��ld��L�hߖfD0I칐g'_v]uy���#��T�&�I�s�1!s�� �F�J��� �Lx,׺�Ơ�ie7��}�`��VݒV%��-}sŞF�~�K��,����ٶ~�w�A����(b�����z�Y�T�S#^�r&�bvۿ��,�H1����.�r޶����z�0������������a�Y;�
�����͋�"d�
^	�x �@'�t6}lp7��(@�YOLup����Q^�0<�s���^�7ӬhU=���v?��W�;��	v���=YG�,ㅃp�I1�d�K\�#y�;�f RB9!����>~�[̙{1\�L#"(���ÆS;0'2�p��<Z�VxU�+r���#���t��*5�����^��{&�(j���JTpd��J&e�]f�zc E�ȧ�<���y9B}�";��|�{�Ɲ�(����t��_��N����|Hȵ�/oN	���bs�������X����� �HB��+����r�����ױ`6[�^B��`����0�#/��%B��Ʉ��lv���p*��/RՍ�d�q���2� /{��lG���'0E�jtn�9J��h{����=K�����5�3��7� �Kh�*aB�bR"�e�����c���4
u�Tp(��r����C&�wW���fF�gQ�$�J��4{��{}�$�!̥f���'����`v�����Ĉ��|�m�\��铄�\~��AK~$��2�ײ
�dm��:lu�� �>5\L?��ц_+�7H�ʢ�e�=�;��F��-�r���ljf��@��',j	�mw��;����-�Gc�O�֫[�<f��j��G%�(�P��	�+S�Y�n:D�=�=:�[`�ι[#fȨ�*)LωΠTDe��V�D��kWzǅ��#$��E"t�f�.P!���-g)2���|	�m��J�ס#Ƶ��Y�Ӌ���`c��q�4؟���������qL����H��~�#1�p�č8�)o�"4.�Tm/�#�)��u �j�c��.�q%��O͕�Ǯ��,_n%�9$U��2�Bă+g;�u���4�oBb�������#qH������$�}��ݒ+�x��>��y�+��k��dh�1�D��R�A"��U>�2�"������T pn�Q�*�	������L�P�ߘ�(++�0��IfF_�*���ۤ�a�۞���%��h�B� S��!��Q~��^ =��*;S0��H�2��s���3CN�_���pp�b�����A��ϡ���%�9��O([��kv.+JL�73\��iT��n|D������s�!H!@0nRQ]a�B�w�U��x����!����~�x�:�H�ҙ�T��V���4	��cU}�D��7,�t�DXC�LMh�y�H��T����أ0)�g����16*q�Abn�	l82�1å�7�)w��ۼ�i>[I��</7S��T"���.�@~O������%יMp�ʡM��Ѿg�,�	����P9l��H<��.U~���e�,D�x6�E��*;��C9��OI1m�!q;���۱p_���a96~4�&=xlP��;+e����j�Ru��g��qN˳c�o�}��ſ�X���Y�l��]-��	3�K�Õ?�C}�e�^_����U6a�����rX��&"��*�(�	�jTV�j�����+�,��԰�h9�
?'@M%{��Î��qdq�D�W���l�U�o��,-ݩ@M����)ٕĄI�5L��/,<���O\mM��	΀��"��������n�g`�4�gȠ!!��)Z�Sv��yGP'3[��5����2�q���X@<"J�z{CT7���k�@�ܙV� ��h2�WWy+����c��w�E��mk:k�˽-9D��6wӥ�dK��y�g*�ջj�s,�90a�0{.�xq�!�c@��S�}�i\�����A�g �x~=d�5�\����Ħ��HS6Ԓ��=��> �Y�륬���:`/��Y
d[�w�t�n'@�$��|�cǁ�mK$���b©�&�Q0�s����0�I� ���!��� GY���}��sP���s��`�t0����H��h�I���s����q��/�{�bUg.z�d��I�c[�/���:��r�@�+�^n"�GzDۧ��8q�� ��Ȗe��N�fB=��'����q}�=�b�'������0%��GI�TX&��'�Q	f�_-ؚ�R���VYlBP �mf5�� �<�{^�D��`3���V[�r$���4�� ��&�MR�ڶ�g�O[�u���X<�&����u	�ɭ�g=��Vo$�2L�Tޢ(?�͘�PÆ��{��x����b�J�ĺ�"��+�RJ- ���p�>�`Tlrqq:}��� ���Cj~���Џk�}z߅���Uv2>��\!�4�]L�C�����^@�,��������� n����ӂ''�
b�Tp �>��a7�8[i�h���a=��r��,6����i�:E��R�(s��؅R�L�vZ��e�פ���?�8��$+'X5"LH؆�5�̖Sc?�gq�Uo�@������ШBQ캴�� �'��R���%{[��m�yujB�^����YN�C �ɔ|$h<[��6�H��#�a"6�k	>H���_�P����R�{]�ou�J���8��΅Gį�Q�����6��c��� &g5]���d�����"�Է�;� G�2-R�gȰ�5� =�z�(��II��3�E#Qč�tLA��_V��o;���$��£_�\��?v�_Kӓ���ѵ5GQ�?�������F�^^Z�H?��Ȣ����� ����~�*
�֝[��qh���͵�Sa��7��
}c�z��z˲�w�����;�M���(��g�+ؙ"�����O��w{͇w'D�epCj;WD�*���X�GoƬ.�`��@i�X�aZ[����w�G�D���|��2x\5]G��[dG��$��t� �w���Q�B^]1� �W���T{�FH����AoD�&�����/1���8����A4e���#�
�}l��8N�XbN�;*Q��v��lb%2�H�����AC�S6�S����@���"̗2?�'ro1	�;��#��S4���=J���r�w�FiF&d����aF� �-�
��RX�$�9�W��$9Š�'���h���`A��7�)��fh�r�b���*	�}�?�?�sZ����`�\Y��^�{��&��	�u]�%�C�S3�;���
��|F�^�ׅ�%�NՖ|��eێ{^<�=����8����s��No�1���p/<&dK
ce�M𡉋�)�ʖ]Y�'�i�?��l~�� �E��7���{l���S��a�V��@����#�%�v>�U7F�dSi�|q�"��0�7�7<�/Ώ�M@�kP�ml���0L��P�ıI=��X��o��~���D�G�?O�S�������{� P���b�w���#����9��`��9͠7D:sD�T�X
�R�N�~q2�I�[�q�֋�Hf�z�V��BY"({�Τ�|�o����N�NU��$:�jؙ�3^m���q�:�Ub�n�����@�1R�N��jҐs�a���(�joќu�K߮�C��&�[�qoK�}��'�N�I�����d��\D:�Te4+B�Qj�n�+5�[���4��L4�/C��Ža'y{���c�0�s7�e�G	�O��d�u��}��N�XOO���A�������_Kz�#0���l^�A�@�^�m|����e�N�y.��eCd	�K���;#y}��V�����u�U��#�!�k$�������A=.Q��x���)ؐ�h�q�p��I�xO����z��d�K�!�g��r�R}�k�r6�e�X�6FV~�����Ӻ��ԲMt������/���,�n�(͝��u(*���S|�J�[�͟�͒.R���~�� l-���K�_6S0~����w�a���j�B$U:���h
g��'S�xix�?��Gw1� ��>�u9���>ע�&��	����K����0�T�)�Zt�� Ҳ�sdt�
k�xdӅo�WA(~�p%�����}�@`4#�cI��	�N0rrqGFz���4\}[�mǅ�5( ��q�GB)�:��̇w��s�>сs]�U���o?��ڼ�L�%�w������k��F����Cg������z��m`"�
<@X�CԶ$b���֘΃��"�_l�u9��w�yuO�:�� ~���pzk���Q�EW�~?�f���)xQ)��u�ţ�q5�z�p�+����U�~�4n).R��y�h܏Ы�����y��ú{b���oX[`g�5��~D�0�c-^�6ӽ�؂��ze�	�V,nac�f���]��$��f���������Ml�ۉ�D��|��y8	�Lh�V��$P"��B�Jv��vK�o��)����Znr��,�6`X�]��$�����mV����b���Qƙ���r_�����N��{h�US��Jo�(2�̨߂.k�{|��#)Q�RV�QZj]��+��(P��.�������7e���68�FSdJ����N2:�`Ͷ���7��á*)$ۍ|��cL��t� %��&�M�v\�@z�#�|�L�*ӵ�-��hNeDms�*��9���ւv0�P�K��������p[��sJx���OF?PD�5��N��vC
bɧ����+�~����dn���8B�]_�0��9C�^���,V!fi��8w�|���S�#~���D'Lrc[�U��(N��Z�oc��9BG(��Mj-ƀG�d�
ԃ�׾8�ϒԽ�H)(J�� �(bb&@t@����E;��:��}����Q"Ŧ�I��&ľM a��+G��ڪr����֫�y�_�?�v����Ɔzf�/G��A݌3�3m��\��TB�t� lr�O�seK���|;ㆤa���ӕ�=̊��9�a��RU�H��Whٛ�x&'����e�8��N��Q�|���W׏&l�C�rب�{,�A�v�E��$�"�EhD�֐�<9��+*���Ž�	g��d_��.޿@ν��8Q��9��)fvǉ��Z�.*1ex�pOB5�x�ʆ�=�ՒZ�����]�~	#�0���k
�b�&�ޱTƋl�db�n%�����faz����q�F.���*�
�KBG{{}6�#x$^.Շ_]���J;��iS��x�F�9.��uX�cl!V�����◮i52�xf��h�ּnXm�lPKl���AK����k�ҳ�YR\pf���ȹa��S�&���H�.78޲��@݉݌f�V"ql�u�� $s�źѤ'�cjd5���R5�$�����W��0�\����r<�|ҢsEҷ��B�H��yJ�����D����v4|��������1�,�x�A�
Ļ�=�������A�͡b��<{�K8��~kPe�	7���X���
9�g�%
K����)���LFk8���֧f��PU�`Ə]�w��u���_�y�_ N�1�d�I'�-t$�"/9\n��w2dWҀ�#5�d9��
*; A~�?�ֽ�a�
���5��ʸ���t�m�nd��	1%ʴ�P��=6E�N�^򛺱���%*�Ag�E��ZZKέ}��P������2�
!@����?��*�5�U���Z����7��³�����S@3*)w,���ᵣ��:��<����tῘ������P  �\-3�#!:�1�X���f�����;8����=�W� H����$�(���^
l'���\@�t�B�{}5��(_��6��m��lg��Uº/9yUpLsW�i}�.0��o;��������㠵Z��/�̨^��W�������} =�5�ԇ�(^�l��= @k��`�F�9泾� ;�����)�TK�Ŏi�)>���5 D\&�N۵����H=#1���d-6�ծ-���'P��d2����W�{����b?�
X�z�3?�+����B��<%�mb�ˊ���@�	��
�G��8����;�9H�M��u�C,��9�#�b�4���`���d�����l't3�DD^g"pwE%����ŝS���^p>�d;-��e�����_��_Mà���U��SU��F���iV�}SeB�)�t#�M��=�;7���P�����"U^���?��}l�h�����̑�ʜ��le�P�Ŭ\����|c}�*z^�)ӷ��SS	�Fs;Id�A���d��w���-�L����4�F¢٠�3��Q���w�6�Ū�]nc; ��(/�W?�n�=j���uW�d�l�T���'���I��Cҗ郱��������{���T�H�[��k�f3iI���&{���Ӄ����!{�����/�'d���ܰQO�#��Bl�V�#C�r�N!�mo�5 ����Z���Պ*�G��v!=���з��ګ���jݖf�^4ǁ�"�(�w�I��9ֻ��f[��+q�j��rm<gq	�f�"A�ͺ�3`Q��Tr;���O2��O�~B�4�]�)E�lI�
/ҕ_Mq֍Y����]@�aۓ���'�ׯ����cv�����x󦨾,�E�\��ɣne�m�<�f-'5�5�yfq����R�\���:��G���O71�
r��ۉ�s��c�n�%�� '��n����A٫�X���8� Uq�o1bՊ���.��f|q�jg�|oU����|�R[:@����ʥ�~���x�$���|�t�J̕���p������g�71�=�J�R���k*�$B.���r GB�㸧�)�堚,�NE2�A���1��9�\�7�ϊE�Xa*�/��4%�Az«��H��>��gn#�K��B΄��z��0I�Zx�U���h�<��=��/���Z��B�`l�l:�ld�1
o�����(�Xz��������%<L�b�jɄ�(�5[}a,?��s8[;a:���-*�MVC��A4���<��8�Z-����
�_;`�̲O�h��@��~�w�.f����)�5heNo5z�at�YϜ�C��sÞ|��
R<���$�l��k��DSE�&���Â������킠�����+�e��p96gmӪv�.E��[�B�l��O����0�Kn����L��鈱��t�f|4J�p�|��Ú�W�p�^u?� ��삈�o�F)��uAq�3/{����hq�7̚jg�xJ������`ѱA8qy�_mY?bS�p�$��bl�9��.�s�<�)�B�<E��5���R�HZ?xD��2���wS���S$p�|�� �yO \%��[p�����Gc��!��_.����u9���=q0�<�
�&*9�'����=��icί�����q���O�o�R� �_i�^FS%�b>�{B� Y
njD�?N2X��뢏/h3M���dRT{W�K�0�'_؇��A��]���J�:�w�7����m�j��l���\�|�v�kC��[.��~��`)��2ut���C����HN����(����Ĥ�Ċ��ϳ}�S�Q��y�"����,��7&3X6�WR� �U[
ݦ�c������-��g���i#�&k0r�̈��/ֺ���3���v�@d߆�asW6j��8j�
g�1P��+�����>l��[v��~�������IbVߧ#U�����)���~{(�
ǂM��@XMP��c� D����z�i�d.�ΐl��5�wu[?�s�@3�$ ^m���_2e7: �p���q.��V=�a�\�يg'1<�(�E��C'�~a� ��T�W�B��sY�];H7���e��o�{W�\����kp�}�6���+0�2^�
�Z��ί�pn̮��h�!�Y'�:�CX^��&?6%��g_�)yՆcݥ��鉤)P8S�n;jW5	��Q�`��5å:�b
X�~�7�s���:`��׺����x�[-����<�΅�����!��Fh[��yt��>7\b��!�Ӆ����@	ơ�ں���J�ᾚ�<�2��R�kU���@4�i��Z��I����ۓw���r̘���p���
��p�P�xh��f��<�O����]�P�k����B�M�=V�J��	ț�Zlޯ&̓��GA�Ӈ�����yч{�M��g�o1řׅ�N�@qf�8bP�*\�[�˵)��=��+ֶ�9k��
�Po��36��jN#X�˅L�T�
�٦�Uo�ڀ���~0�����=�(ű�O|�tN0��y����ؾQue=b�egq��?�꬧t5���W��T5��;�d
Z�K��+�}��(��ܿ4�ź=t�_����%"������f�J!�.�Ϋ��b�K����?�A��9�4�ZK'�
`^�0�О�{�׶9Y�)2t��M�^���̇@���6y$�Co��ѳ*�_���3����:Ы��	1�6jE"�R�c=�����=%TJ�<�<)7�cQ5y�ߎ!��V�v<����Y=�>&��� �Y	b+ � J��e`H2��jFJ�2}|��\���4���[������,����x{�>�
���Q���x�F&w�-���E�ݒ����o�8bݕ5�\䕶ޅ6է6=�%T��\q� �I:�|�w���I$r�z��g��Q��֘(p�n�An'++�������UZɚx�?�
�y���b�2�tQQ('v,O�T\�N��j҄�	�$���8������;@�;9L�
9����a,���fe��r{]�9d ]��S+AC�N/��vc.ւfya�������Jm���7�k���yƆG���b�4��������ɚj11�ɟe��_m�0���J.f�E��dWBH}��;�ى���i��6��\>����H��@ұJsFd�6�����S����s���
)�k�#϶���mA��#���xk�t��.��A����1������ ��u�D�_���d�]�C7]#����:y6I��+=dqs���z�v�o�d= /EQ��yL!h�1|���*����Sv�S��F;"�-���W���Qū��g���A�|�$��nV�Љ����Z@;R&b`A�=߾��
�q"X6��5b~P�c����*b���O<ڷ?��n���8����� w�x��M_����H*:��i�)�r�b�ʽ�����h����R�u;Hm�pЛj�Q %��.y~��-1�����:U��`�O?i$}��Uw�AA�\u�%Bۍ��A J�,�DB8C���g��k����Rk,4vgN��r�Z��������i>�+����-��[�!g@%�S?bC�sA�ݮ��0�i8��6u�ր25{�M�2x�� k����q�b1q`���.g��Y�����~A��E�."��t^ȳr�� ��M<�qn"���{�����Xـ�l����,lP�y�{��8�5������K$��=_1߼�&:��G�GL� 9���{xj/�
Jª�D�2�/6���!v2�r �`]��F��S*{��3}�ɐ�y���'ǯj��a/�ekqW=�o��}�� �c"ΓĴ��1�g:~e�騕a��|�BͬC�9K�g�;�:����	�<E��\sW<N�t2M�3y��bM$��t�|qo(!������1 	^���f5�u�cbm7Ɏ\��s>}O��6h$(�W�[�I�#4��2|Ƣ���w��8������E݈*�#(��E����(���O�#��&��S"��qe{�g^�<����P�}���=o�+��Q�
hZ��k ��&��P��ғj=�gN����{ç�|�w�s��Q!L!�w��kn�cV?�T|u&�C����ke͇�����0S�XΎ���� �c@�4���=5}����̛�6==�Td�6z.�טa��F��ۿun^A����.\�� ��EPy�𣉷jq�8��~M�����j V�.��hS� q���-Y��'���d����P����~d�sv�W�}yfU�������*~>V����Q.�-�3j����jH�Te��u��~���IԀ��@huɧ��*McTqw��,MEB�f�:	��0��$��t�e��9�}��S2p�y_��_&�����i�AoB���d�]�+q4p�k�Ys���������[bb�:s��FrFs���SIP�Ҹ�;�0�7�R�	P�6(��I�E�+?d����y� m�K�'�>`i�e�v#��e�x,u��-����{LXNRϵ�o���p��L�'�'+󑖽��`7  ��Y8���3e���弓&���ˀ����ǲ���O��v'��a�������Q�*���-��̑Ž�:����@4w:�OY����j-̀]��*y�߮���M�M��=�����jD�TEP*%]����̺�Dq���|�Q��=?FC8j���A�'�a���KN��ң���h��A��(��>��G|��z<ݤ�|���~/�3s�Wv��O ��;�ƀV5����[�O�[g���vuc
����O-��*�k�ɝ$ĕ���<T�y�%VE���h�|��>�ÖV䴽;/w���Ŋ�թ��������j��P�PR�r:~�+xJ�t$�-=1����9�(���g�ѐ��CW!��!����!#L��^0�kؚU�e���J�>�7���Fng|��YJř-@�3�`���L�(�"�����B`��Xn״����w~XQ��g��Q�ek` ঀ����=́՝,���'�=�r.����v"L�Wh�B�7f��R���J�!� ġ�@B�6Ԃ�M�9�}sda	�R̹�ɼ� ��0�-��Ǔ��տu:4jV����xeT������V�EQ���s�@P�t9Ğ�Nٴ���K|���U3��{fW^�aS���^;��� w��ԝŝ{����Ρ"��p��L���iX��ͱ���_��쪀E����`�
@bB�{�x�_ ��7}��5+�G����,C�L1<ҥ#P�(��I)a�,�-�1�Ez7A���3���Aiv�o���A*�mҟ���6�?�L��^�iT�s�]���c<^�Sv�!J�J�Zp!����I��}IN�.�ǯ9�F��9ZZ}_���<��c�в.�%n��3����2�4�V��n�G�Q�͏>+f�FE��q/�~)/���iH�s"z� �s�Ŋ`��;��J(!���B՜��.P�g9}�4=j/�*��!�=�����	���ǆnS�n[�^��ը��]���5^�x��Q�A^ԣ�5m�G4Q��=#�m�)n�w�kU���<��Mך6ペܐg��� ����ɒf���'��A.�_�s�u+��+��*JЭ���ǡ���8��&e�w[�d��>4����e�I�jz�>��gL�}�՜��ǖ5\���_c�hk���"���Y4�HVz}��Q���b7���?�ڂ�����щ��uGg��ʺ 	�iz*4��(}ֻ���^�����~e���I� 3,b �wSnO�E(c�=��P%���r�j�6����Z?];"�fhZ�[u*ZL��%e�.�5��k�,�=yA�}Y��
Y���U{U�_^PmO6G�W���l�P�Ie�33�ݏZ፜~&���"��R�n+�-�1�?>$���a��]��Q$��1T��z���#'��J@Xk?����6�P*�=Dᔙ:�"���(�7%aqUpw��)����@�
����W��)�3��tm̉z� 	4,lVq�H��AEi����������M�<�uޤ>�5�cq~  �j�-���7�3�2X�v4���M�V�x B-�h�B�����t��W!���Di�eH�b�/��b�p��b����`�d�"�%!b�R������ܮ֒��}V���4��j��c{�8�rWG�.=��e�\/ٱ1"��^="#�}���������kNBi�m�H���n���<nr�1�KN��@ws5fR�)�%�{oS@���,#��{(����j�?̂�o��>�k3p�=�D�Ux0��+��K�'�2�W�-g��k�	�TQ��J��'SΙ�zM�gk2Y٦7=���c�ci.������q�PմG{��&�+�� ��N���!i�6��4(4��k��N*��Z�{��v'���p�)�e�b����`]3������	x��*h���]�<��C�a���#��(��X�$'%���#$����Թ2��!3X�g�p��{�S���TA���B��*ݹ̽d�aG]$ ��5K�H��_ {�`�c���a����>�](��)#E� ���NC��ax��/�}Ⱪ���"L��}�򛄓Of �"&N}@m,6�4l]�8y��XT�S���+��� ��V��́M��5��:�o�{��#�+GYe2�k�.�A �YZU(?���U�ã�'��'~�R
{t��^�S �B;I��J����R%9����j�.2<�	F6/����ƶAau�*?0(Ė���&���$���xO�9��q���Ī)�'�za	�tۓ~Q�!�Jzj��W���#�Ё,��$�7�d��
z��|�J}f%���'5T��9��/F��H+��5*����[HIC7��p�3�3�l�� 6��.��f]�]��,�w��+�b�q/��t�λ�P:��Pr���D���A����s(c}�R��_T�\w��i���-s���t�Du��h���e���S�n�amg�L⦕(@ �古A�\�s�?ۢ�m/?L49&'�tl�C�)�V��x������Cc�N}��?	�sA�|�s���T���=��R��q���v\��]n^k�[O�o���@�A�	4�������/��Y١�񝜚�g�*���xFL{uU.��4-��`̕�i]��.{tH<:��.SH��S���ruV�֕�ˣ1�)ޟ����7��&,�.�
�+�:�]�ѹ:j"�L��%�v�k��Jh�&8[6%e��j�:��}C:�^f�Qv��Pp�"���-���v���$�H�,S��/�LB\o�@� �V���,�gR��Q��`E����e��Y��_1v��GuU�r������p�������Ư�K%	�m��eS�TBEE�R���TN�����^3Э^6f�\/[�zc��71��,	�g��SaNB�[��}ϴ*j��"h�#TI<;<�����/Ċ�oQ�xB�B�T^��E+]pl�tx��H�x��U�ɛ!���<�X��?ý��"�|���6u0=Pspa�g����%]�fȩ�-��Y����N �iW$�D��*.��!#�������R�O8XsZ����ِ[�s�_�'��Y�*���CsdY{쌳c�י��G��[-����&ԝc�9���?H��RD*%��m��p�]!j��28��v�/$nRl��@[�X�:&��U�Z�(����'p�.��rA�Y�� 'ȗ���`�CU�bB�
Ւ�w�Z7�j�-0��X�����>.����p�[�:���Fuz����g�\����H�w=P�JTTα�	=I�o�����O��U� u/K�&���V}8 ��c��+�6�o��nw����S�+�|x��`��_^��	4�q��)J�5rA��H]?�XzϢ�"$��JX��O�EL�AN�����1��ɇ;t���`ǵ�����s����?̏�zl��&��� lm��a�Јe�a��^�a)V�X�O{:��YL�JY�SP}�UU�{��"��u��N���ת5cm�d��B޳��>w_&����^��~�������=,H�.�,��7�grh�HOU����]���B��G�U�[�b9����{����WW����ⓐ-}"�5��Gz
�o7(|{M[�!�sc�b��q2�]���a�t�LA���-�7_v�Z��8:^Ҕ���}�r�	�����ID��U��,j�4�b�Ħ Nl��]Ucx�j޻��#�?�����J.�X_&K��y�s`��"�#
y�X��y�Ŏ�N�^5ޠ"����6ƪ�E;X�(����z�I�l��l}��Z��S��1����5����N>�t!������Ȋ���Z[�uv"�������]�.�`�I����*�g����Ksp$������u�h��ˋ�o�p�Wbj�XrB��;']7�/3��1&4��x%p�:�������<,`�lvs[V$M�3k![������L%��������P�*O�x���Іz�Αyߐ:S����s��X�~Y�.W�?c�}��;w\|�\��VҾ�.17<� �@ht��"$�W��*0��_	P��x5�sñ��Žs2�&唭>�x�������2H�Yô8��V�~�2��.t�����A ,�;��А�ยz��%$��rǨ��R��.q��<��ti�bdٽ�H�:�U%	Ȑ�\z�ii4˒��S*)�����+u�ÿ�K��/�,�����#�(5f�T�eM-|��|��Wpi-��� �*���B�GW2�F��1�͕�/�Z����*_l_�=J���bǨ�O�\�	dA%,e�1�D��c��$j���5���c����X��J�B�ZpE9�W���z?�����Ꟁ@��F?��z�ߎcGɰ�	��B6=aUf\j\?�)^�<NX1�qCR�W���͋���#"0N����~�y����rm���"K���;�d˭��cB�\8У���Y�%�R�T�:�u���ڷ��q/��2�H�D�0�$z�\��h
K��Y�*:�GMX��n?�RnKc+�Sڪ��hOmW�E�_�r��N�V�ڶ�"A�.=u6�w��6n�΁�M��h��ȍ��<M����ڻ?TQ�V�;d�O���mܖY��ɹ#)>t�\~��ƴW%���?0<4#4��^#��
I��HԴ�@��Dڈz���ON�P�3�)b��yZ!�#�.&B̳�eU38[�Weȝ����g����x=��ڱ˓�3�:���]N��m�[�a}c;j=��I�ʎd�K�.�5��G�^�fyc,����2��-9�o��������.�TmEo���
yo��Z�U��Z�oC�����^D?4��Fw�U�e>��m�����],1�/���p��D�d�N�ɣ�-�.�������Y�Egq/�GSp>�72E�V�/�X*���ɹa����R���R֌��M�T�Y��8�����P�\|b�4��9/2�ض"]t��V߿������n�q+7�>(f��T��)`⿄Jb�.���v��\d�Ldo(�*��f^����yH�鈍K��)�:������S���fM趃�u�?s	x�����qm�_s p`2d"�d�
�V)oaoU%|r�>��y{�o��S��1�+i�&'��R!�h��K�f����Ǘ��} ǘ\	=E�����[�w�d|�"�_�����p��d��֖�}��� �*�0*`r"��4c,2��g��1r�L*��?{���Ԕ�v��=N���	����U���EW쐡W�S)��1���T�������3V��c0�i��+���a�M�Z����z���a���b�*m%|L�&��ЩO�}��Z�{���=���|n.���iq�ζ4�K"�5^��/��l��RmnDTOF���b-�n[�����V�R5PMq,ݣ���D3r�����>��0Q8��$��ݦx�k;���*�I̱�
����8L:���=��Α���v	�˂5��k��SHZ�FuW���,��v 4����GI(ZM��
,L�03�͕%���m/����zx,��d�o��~\�����	���I�O�T�?K�`/rd��LMT(H}��V���(����������>�	�G��OaxC�K�lTlR~p�8��6R��T��@l�����z�Jj�H0��j�G��5�yB��z��n#U�C0�� ���ԅ�B��id��e�鰄"IZP��ڊDn�������&��n����q(iX�M?�Mq� _R�"�p�D2@ja�~����m�~�-H����]��er	�f�,���N*zй���b���	���Cu��l^b�<����D3�Aвr�d����ync]3�C�v�2՚��K��N7��	ܡ��dh��nCCTإ��.�+�tB�n~�:é��(��~t���f��$xF����|�8�ޙ0�|ۤY0od8oҢ�dF�΅�3n���ޓg��C�yX�j����F���d��*����P�=����0b�~��7Ƀ�� �R�8�Ң���,���]2���~{�����1�	�EH1m�"r�gUn7�	��k|sN��o\�ȶ��t��r�H�W��*����q��."$�?$4s�p��~a��f4�gŮ���Ą4�br2�?&�i�ۧM$_+w!!�,����46�W9J����}$i��:=�w��1���F_Y�#c���\���Gi0:��rJГ���Smd��##�"aʲ�����{ⶲ�S����i�`�t(ϹDl\�IC,n��e4%(߹7y�c���U���o|v�s˶�tG��@i�� ��,��)y����W�|V�?X��/���"e�{�U
uN��&	 ޡ)���`�)�v��e$�Ad��`k��p�8K��p1�� ��6�z��:�L)�3i���q�>N[��MOX	z��5~1�y�޽��?Ϲ3P��pAQ�7H��W$�_���5(~y(��f�8�e���=p�ӳ���G�I�iG��X�^E:���Y齘��G�2K(W=��p�M�p|�w+� ��;.,�$
W���Xbz�I�|0�$�$��z�9Gw�#=iLru"�W�W�*�������;H7�=I>�Q�!��a�©��T��JQ�HI���](ٳ�'�uVhgD��^��C�� |��;��$_�X���?SK1���#K^Όv�_1v��jt+n�h�MAC�iX|�YxE��Ͱ���U�aǔ7��h�*?�*�A�rXG5\~�6�*�����U(Y�E|`�3ߢ>톊�A���T��1
1y�#���YǕ��3�{d=�5R=�^���u�2�����9i�:=�ym�+Kb�q�7"��Li�����s��@��FU�o�O���A���}*n��'�E���I���i$���~V��M��G"b�K������Q��S������۔4!���D�e|2;�|:�H�g��c{}R�zw��Q_''n�_�]����l�L5�7�ۇ �/�[�Ft�9�0'���ج�� ඈy����%5���|�O�q1�_v�!b̥�(z���'�hg�<�="����H\�̊�H�mB�P��w��!��q�>���?PV��\w�]Ԗв(y#�m~V��gS��?q�\���$Mqe�_c��6���gEEw�&������7>-�}�?򵑰�c��r�H���V�c�3J�_k��j>N����o���5��J�����M�`��M8eZ�2��]U������`DS��*P���5��j���Cf;�O	y���x��iI�@!�D��]�V��ß?������ʾCPWoxg�::J%K�:D�1b�7rŲ#y(���u�@�I*��;�IOW�a�#.�u&MY}�P��'m-��s��B& ��d�e���'�33�2�Q������z�I�	�nT�8��߶�u�<K����.M�A����x�s���Q��q�x8i�����J��p.Q�.��h^�Rw9�kP�U�����68@[@�0[�1�\O���NK|k2�>��<9_����]�M�����f'���p N�k��j����˙H�i��ŻQyڂ�[ʘE���v�gG05k9Y	������
W@VHu��g� ����!Á���⻻A%��f�����|j?.G�����RD� �J�;�쪱�L��7[�'�s���������+��������d�i���k��!t �h)t����e��J������&��'�&�ZH*(�J����&�˔OQT���~�WH�aܪP�U���P#�m���q�P���uK�?I(D/V ��e����C��"·t;��+�*W�}�_���LE�������%�?K�`�I�ß���^2dn�A30P�=��WLtL��jE@^73u��W��_(����ݮP�<�ɿ��hyQ���:6 �e���Xt�6P��s�2�&�1  �z�XY2[W���[~�Y�ۭw�1���\�Yْ*�%r{o=�P3n$]�u-E������a������y�ȥ�c���L{y&�y��w��⠷;�Vv̍so>��5^Oc��Wx�zt�Gk�)ñ��ޤ�p�7b�]����^�D1ٽ*L��BA���z �o���%n:>�(C�*S�1Kw��q�jFh�ɐ���K�sgr�vT�yآu;0/y\7D[�|�Y�3Eyy$���'ҷ=�m��-{}�o��Ԙ���$*5�7g7T)�u�ط[��'�Ֆa�U?���8XBn45�L��;+�SxR4���e#H.�m�3�08�F��9:���П�1�$�Ȫ4�".��G3Rs�o�<�{շ:�:8��B�5�l�b�(�.4�B�.�{6�u���-^mÞ>�}��܁��y��A�Y>|.-���$?�s�7�9�(�m� 1�鉺YF޴�ՠ3��w}�����|�X��x^�$��A��O&�g������| ~�+�E�(�L.ǀ%��c&�6�P��Oz��D����Lc-�1�@��e9"Q@rށ����;�qM���j8�W<w�$"����wP�8�CfI1.�]DZ�4)�g���!�TXV]�?*�R��"����$~T���G������I�Ct��q@�OHh��tN����%���ﭰ�4YC�ug�GE(D^b��\@<3�آi�/�ʻ����4����k�3��DG����)���8�+��� ��E ?HP3��f�5!z�'�7�kX�]5�/6%�B�T���gC$i�? �\/.�>�f��`J||�ڴ��p �x/0�ޘ����̈�.�f+�VF�._T���7����'k��u��^i36ØN�s�Szg �ȴ����W��T���&Bk����N����㨮�dd?�6j/� G���Ҏ���(�(��:���D�0�� �ȰhW���KW�����K�F�]�PA�"q[ɻą��$�(����F<d��3����3��z�u�Qm��f�}�ܕ1R/����}ֿ�u � ��������6��;o�g�%l���y����	f��O=U�&��T��`f�$�	x��*�ޚLWU��q8M��s5��K=�C!X���o!�����o�?�|0d�A����:�۟l@@�/:��Uq"A>Nw!�&�Z�9�sK����Ǳ�:��85t���P��徴�1�
�m�(ڥ=��&h������>Ul,R�\�:	0=i�Vh�c��y�;�o72�߿}L�sD�d�gmw��,I�����ř�[�<����L����:�$�gaw�d?�z�_��=������D}�w��;2x0�=��Y-���c�&��5\�M^  �tk�x0&1UO��g]��N�#a�w<���͛ R֩��x��Ed�یu��w��5<l�U��qȿ*4Y���-~D9|��i���}�iR`��0Zi���p����{�d]��j�&z;��tO���U�F����$:�_�j���h}$N�ST\�z$�G|3�M��(�q�ΰ�v�[Y���u�,�w�E���i
���1
{��ڊ%in����z!�Y<6	^$����F�oe��۳5�� ?.pBi����@��E�bU�>ޢ��U��5r����{w�����
����,t~���X]�_��ڥ(�d���6����� ģ�=@�&��$ �bS�c���E��O��W��e�X���<\�������f�A��4���P}O�Y�s5o�
4E�@�	������1��'Јr&Y��D?z��@���,�t���7g�!ԣ��(�+lC�<��Q���h�=U+~^j5������a <+w~�3��D�'-3�zc{^o&ȥ��*ݟ"o�J�~��h���
g~:6�*8�����q�#s(�L9o3�x��v�)/q�3�<���g�Q�	<�+��e��Eӭ�H*`t���Ʌ3+`f�,F%���A�G)ȑ��+S[���&xOQ �e��QJ�M���t$¶S}u����l�,�s�-����j��R
D���N����B��o~I�ۯ:�a���<_*�/N��,��|;=QQ��������#�$�8�. �>/��j�� 
0�9��A��6�f��9��8٤�H'D�pE��������E��sҨ�B�u��]OPR�R��We=t�����{|<V:�à��Z���yjq��� �v5	:�r�������ڨu�������-��@���_�Y�8�Tv�)��w��TZx�������%�-jj��GJ��XO�ZZ�t����R�Phͯ��[���u͊��+T���S��e���EB�%���rhϢ31���*@�ލ���w�t�꣞� �/���"�G(�^����cY�7�����[4B_4�}��J�v�Cߤ�z,���u�Mπ��-oCBL�<3�O`�T0��v��d��rb��gb��}�<�P���_W�\��Ò��FOBWvI/�$ [�m�wu�V�� ;2��>+7��םzu�w�L@�6�ì�v'l��̑��cUC	����y�����_)�F����?�H�Ɋ��t����6C�~P�A�1he�,��r�b^��m�H�o_4O�4�HX/F�.�-��E�&I���Jܺ>����)N�-^�v��»��v�ař���?<�{)<�fSK���O����y1�aw.;��7�:���xl�bv`�~��,P��ʘ�y�2�����	4@�$xpl���4��yB�gΡ(�v1����Ɣ@��|��w���{Sf�����%���z�8��1��YT[�D�J'(��`<�64�����1�+6j{�B9�	�gt��D/a��������S�oenқ[�	����j�$܃���m&��U�4�89iR�:s|��d2$5I�1�a���F*�6�`�r���t�?�mbJ�H ��au]Ib��8���(u��Ʌ7���v�n2c^�C�L��=�HU�W6-j�t���	��Q��\!�`̧ݾI��+[9fةLe�$Y�XW�S��MRd&i�}��s)ـ���TnW�6��o�O|�HPڽ�wQ�+���:�Cb7��1	�\1G�K�(�q*�e{7����*Rf�cwWv�Dѫ�����"j|�n8�w�g��w�����Ef7$R�Tio�	�M��a۰��)f��P�Ӑp!e��%9���v��]z���ƽ�&�ܴ�{Rm��J����C-M��y��/��Ar ���|�#�:�|�=oݞ�D� �V�:����G�ף��˷՗�i�6�K��U�WI�_A�[��BL)`҇$����cT\��p =h�|_�\D�BaE1=?�x��_,%�h��g<�z�s+1�)��Uي��� �*,������0�b�l�}�Gѩ=[i�U��m�����3o4�N�`[�A0 �_�h�0`[��L�>��Q�;k�ĸ�*���f�����{�q����!y�3���d��L��yg2j��'|���gS�����Bj����E��{'6���K�x��\A��3pDvh����l �Iy��������*��L�đ�R��aܽ̅��6y���(�'!#�FH�$�r*�N>�x�IP�(��Dt� V����zM���iq�<��R �]��3�Y�d�d3�����p_�'`�h���C#t���%��\���q����na����h���	���Pw1��5���=����9���oo� Y���;�L�Rh�l�s4z�@SfL� � _�����;)�h+�\������ܲ�\��!2L���0!a-2r���z`����Z��X�U�'�Wo��z���s[�!�����^Nþ���-����(nU,h��`����1�A��"ţ�>�ƾ��.pL{�����Y�A9�S<9�>�{�1qf&�th�N�m� ^��u����'v��)�2��Yg1���{�f�ǭ�i�y�p�WI�.ρ�A|��R��Q���ak�L�O���mĻ�#�����?_�S6�R\�S1�b�ja�FQ`����Jp

o��/�u�� :팥p8S2�u��7�5d�E������uq��X�q��$#�X����jF����0{ݐ�y�m�:	���Kհ&"*���Vo\-Q"�+�Է}|X����_���H+P��!����(�3D̚Hc�H�����@ʢ�� iD���sQ]v4ڗ3<�"�����o7j�M�2��3Ħ|1ګ�
%����G�@u*���K!F��]�)�A�M�	�����ݷ�.F�Q��������'V��/����O!����G*ͯd�ͩ�x�8/�}v�J��8��(3�ja��Uڤ�` ���1I��y���ik����.��jl�V�~%��@A�+љr�,@��t��:I��"a)>����c��ƈ��5i@\��ΩT67���G�o���\t���Kžչ�$��.�*�y.]���j*ߖG�!};�'�L����5���������3a���*��?�6�8v=�|{9a�Wkr��� E.�02�(�2ŒE�e�𣙠'd3�7�+\+#f%���T��{L��M�y��o&�x�ĵ�H�J�c� ~����½���ymι�D�Hw�N�1H��gf04챸�����ʡ�DXI[ �����k*RN�Y�`�±=0�o���,�,!3�d���p�!�3�ǃ�w�����%'��7�KCD?��!���X�Bi]���>�Um.�Μ+�)<7~I�A�Z<��F%�/-��bA�=���u-�y�}>sv����X
�D�{���{�Z�&+��0�N��9�!H��y�?>���|%�5��E�tG]�P�D+8W5-m�1DZ�)�2�����S�h�-�(��X���so�d��1H�R$QIO{~��_�߶�.U�~A�A��6\��$�X+sN0j	y�݁Cj���z�V�F�ahhJ�e?o�`�T�V�T/ rwH��/��Af �9�+ik\/0�����)��#-
�8vZ�ws���"� 83�/����K|�_(����B�l㏎U�[{.0E+�v��ڇ��U]�wl,��IHfE���}���݉��Sze��e�����'$�}�0Ledx�hJ�s>=�\"Kg��r���c7%�z��
�I�}��V��b�f����w��5ϾF
�^R��H5(� �5�1���0�>�����M�JY#�O�%83���7�7L���F�.�󥽌��� ���g���m�q�MC�\n��Չr�j��k�9if;��WJm'��Z^�Q��	��cꑼ��*3�Y�# ߍk?W����S����!���]�T{�#s�0��T��TȈr��Rnt���'��!��%�zʍ�dE�^�����j
�Zp�wQ����ӻ��(�?��A����.\1�V��Rٱz�+��@��H�����Do�<p������Е���|�wvaO��C\�$�Q�O�Ɗ$5tR�O��'b�f/��
X����8�R#cftr����>������p�^���c1�]�5�������¿Qda�
Iװ����0 j�=Q�_�m���tyc���x
�,<�Yqb?�`�k�A� =G�9�Nl�+vS�f��{M��d3�9�l���-�4����mPH�o�1:¦�]�b�|�sH��9#��2�L�k0B���Vo���8{�I��q�;��g͋5�mMO�M�;�~���`ŕfc����hߥ��O���x2����Ip�`�K�q���j	My���ڇ�-�-��<�Ґy�(V�d7�4�\�/D�����k$Ky>6�k?�`���B��6Y�mAC����\�v��0�8Z�<��uY��Yw.�c��]�T�)}\�� �*R�ff������k� �<�0�*�?��4w;���� ��i:�-L���/�6��A|�/i�vX�\������hMs��K-S5�Ւ�|��O>�O��\���˱������I\�x�Ѯ���'!�=K?��\E�J�$$"��︇H�\{򛓮�	�,��{�7� �t�A/O{�Q琶g�/��^^&-�3�~���G�2h4��y��/���%t�w�m�z[��7w���
�2�X$�e�7g�����}xn�!���xk��7U���!�R����TМ8p�?��8�������K�eÒH).fJ���)!�Q)�r=ɛ�6 y4��~��A���Y,"進�,�,U�ikX�+��BB#���љ�Cg���~�	o�`t������߼�}�G�&��x]+�"�i6���\�٠ʙ���kWN��,��*��Nܻ��!�����<�1�C8�M���1��K�A�m�Hֳ�u&�O�k��"����ܛ<��>9ը+�Ф�fF�%���Q�dG��6M�?գ!�4+��2[m�z\�%�h�i)'?�:���|�����p�$��x5��}T���ZKz�+Q���zY|���{�������,�-��Zi��ë�N�9X��\R���*�V�!ӵ���Ш���D�dZ�/���_���&�&�ʌM*TQ���� ��
M�?�\�
I�[��*�u)� �;�bH/�{���A����km`����w�^����������=\i�ԄZ\���t8�P�'u�dW�W��H7A�c�t/�j:�}Ж����ƈ;4�c"�L�dٸ?�`z9��%H_7�pq��w�0�~�Z���7�C�@�����pt�g8U��a���}x#DčK�"�����9+�L}0���v��mp-�k�U	��=?S<־�̸�W���Ilj��޿��B��h�5�*yC�[��ͤ�����H�~m���������>^ܸ2O��"�嶞[s��7��o)lu��,�P�,��G�ჭR��D�S�V�p�7��+f�^���kd-�/z�3��Z��J����0rTH�[��|�u��~?�(�~��Y�9J(|k���Zڔr��	�L̪�����S����i?��1����#�0�{���.Nڛ;O���g"��))/��c����H�C�?/))}=����.��΢Y�u2�c��Ɍ�7�X�BjO��a�񵺃��nR��.Bw/�̟�L�Q_�Y��W�H��r0�4�(���uV%��o�#ș��a?�{���ct179�օO>ߴ�M�3f�^��QH�]�8�;.!�C��[�:Z�@�Iu�W�%�Y4W�9
��;3�n*> x�]*^�`����$�N���})&6�/,u���(�}P��C�EЊ�'�~�"�X�+k?���w���;�z�#%�*j����d�����M5$\�ru����#����^��N�B�/y�-��*.(Iq�/�a��t+5_�K�U����R*���N-(ET����ϔ�_f2Ԓ�/J)Å�ca���}W'z[�l�+N硸޽SmF�#8&EY8�>�m�k|6tn�QX�'���_�Է/�-�L�{ 6�/WM���Ly}�xG8��U������I��^.�f�`��i�w�kKUփS+���g4.9b �l�(P^�5Gb������86�ҟ[7���bF'��^���鞗���3���ȷ�_��`����.
G�9�2�Qg�K������jr��ax��X>�u�n�H�o��.	A������^�YH�9i��y��@i���;�l����Ϣճ
]�M�$��]�����[��S�d$!V�RxOY��x�4�+�M�E_Ky�T�sK�f��s����-Zj4�v�z#'��	Rb�0��O��:� P�d���̋�*@wO]�<��5���(�+m_g >imp��'t�I�1�1p<�e<Gg�
�]ܐL�ٙ#��T��;I���>�R_,ս�����0�0�W���.~(�X�(Jȼ����\�`h��Op�ǭwp'���Bl�nIP�C��N�~�I=	���K�o=d;���mx�JZ��cG%5<^ ������<V<�IE���fG��]�m��c� Q�l�9�?~_R!��m�-�6� \Oh�xFh�&/Ea�]�`�^�Lq���x%�^B�k`V5m5�c�����`��%p�-O�M� b:k'�3��@i�Ju�F�)+xl+�A���鬯�
�s��Y-|��V1�y���OӀ�~:�t��ъ��d|Y�Ɋհ������g�c.W��b�j��8s+H�/�Q�<����ǐ(�B7�Xl�<�])0���5��2��I`�?k�%���sQ7*�7��f^,wR�i.O8�&�hlgfB�؉�B���Ј�b�7��-��2�_K�i;*�d���[��,�D�������1*L*�����T��̪�N�tV�����Y��,$5����ZyW������U6������O���\�lMά�{ Wgp�bރŴ�\��\x6��U,)����z)Rr�?+��F4ٔ���R�|��/�'ِ���٘�c�����r��VZ�����t�\�����W����ϴ��������o��c1����=��3���'�e`,�IT~G���^�/�E�je)�|�CeX:?�
E�-�?��pS�@d��K�
�~g�x/:�F�Ww�����=�>h�ͥ��#�H�w�}����Q���K��5Z;�& �q􎿭)I;��#P�u%��S���ɎW[=��|С%�kd���U�m�:���8���JB�L��@�W�gO�����9%���-�.���R�(�@ӂ�7E���qp�:9�U�6�畽:l@31+|�"� ���`�ԴMt�U[ ��5*����`d/	&n�PT[P��&	�u�Z��ǵHe�Qw;�v�d��i��hf�gb|�2�I�x�s�%�T' }l�6��R���Q[o%'s~��642q���s�C�]��Ԉ ��8�זC�@��`&��Ӊ���l�?�>_�|�P�0�$��qAq��5'�q�A�R}�ra�\]駿�,v�ޓ�+����FP5
[�exzzz�u�[�8\S�d�"�݈�3�k]}7|��x�xI���_� ����	�2!�*%ǣn0��;c���~=��],Z%V;�����h`��*�&�&p̯���� 6�ǡ8��*�v��r���Y+G�����6�6�/��s����"y�t#a�ڻ���]{d ]�ƌ]J�4%5U���&��=_!���8�/d��t<��"E�@��6a������f}>~L-�=⭚�/�Z�j�0~��@!1%b�;q	VGs:�6���.��=��d��b����S��޵x �*���wV�LIc�H^X��X��w�o��q�=HZIϸ��Ol���M���~XA9�߹u��WK=^BIo|԰Qm�
`�-5O7�����0��$'��3 g��]�N�X\��+��&�$p<vU�Z��^*�T�!�8��u��8��G�P�Yo����XϯmM���ҽr��,����^�E�F�s����Z����w�N����I���֣G#V�3�R�|�uN���iY��U�2�e��,>�������V0��A���h@\��M2i��!�lҁ#cm*��_3��5Qi���PÑF[�u69aK�{5�����b���'���m�����J_�W�iXjFm _b'�Q��#&�='$��bV	g����3�s�\W �5��`TJ��H�}/'1�'r��2ܺM|�������9�%� �}�u�j�⊠�\$/�F�-z��/8�I1b������K��-�+2�a���K�J+��4�!�Z�ٰ�j���ү���*����X�It���30ԇ��Z���棺M��VC��ͨ"�n�,|;�F�������m��@WP�"��q�����#.
%��nqH/0� ��_�W��tDA�VL 2��/N���T�)��2���Mr�����q7~f��o�}��� �����wuF�c*Q�fU֖��I��7DqҘ�fޢշ�s��Qy) �9���%u�hby@Ų�	ʪ�	��^o�������v�6�����8���4"e�$�]G>��{r��QBg;�}*�.���yq��(��Q��ϝx�u�X�iz���	|������mAz���&0F���f�D[�K���LĦ�cт��bs�g�I)*n��e�@eM�qc�m�x�j��:��T��p �|˰�;��ƯƚDy$�K�Ƶ����k���JN�m��M^y_����i+ �52N���2�[�lS�6=�U��LNb3�=��T�c+�~Ē{^h�,�,)m3F5n�8aX�!�UyPZ�`�nC�s^������ȲumX���n2�p�&�x���h��T�t{�rN-!�i�[����2�"�mT�w�^��M�JP.J���w�Z3��ҡ�.�7pn�ǰ���@.=�.�ˏM�%�炛䋁v��#Єn7��]��[���E�Ou�x�|G��WAQ7-�i�ʦU�/8u�O���~OT�3�b�/��mg�)Mܩ(��`Ж����:��t���2dsX$��b�|3�Q���ay9�{:��`^2*�q���n.�� �/��@b� ��y��n�Vכ�d?���^@Fwֹ͜��ۧ����i�	��$��d��u���o}t�Y�A~V�(�B���m�N��P?��s\:�yܩ${�@vN�^��ɵ���;�f1��z��8��.��I,N&��١>;~3̝N��6̭��]�����=�\+� U�ꬸFսNb1�����r����KTv��'�S7��+����=�3&�ꍡ��U���G��-���,���m��,n/���NYa�$�r���l�u�|}	L�{uy�`C��
5(�yp���G�vJ�i�2OB6��p��F��y�<�i/��bL��d������9;6.���H\	�p���m�V��F�$�D�������.�/�R���K;w�K���EDHQe���ܞܥiX���dƨ�a�q����17���(�=��+j������AʈS�گ쑿�}j{�a�!S�:
M/���H�
�)F���y���~B�k���%��=�����I��:ť߅�X-���ٿ�81��ӿ�[$���{ţ}�k5&���Þ%�������%�Pt�|�l|8Ju63[�ׇ����/>G�#�G��Zn\���OB<�g�`�-	���N�|Q^ǥ����f���:�ᕹ���35e��\��	ԍ,��M���\Z\�6]����nm�)dT�Y3�"#}���p�q�"�[�݌��r mk3�|ZV�܈����}�0���kA#��D�����@	�����PSwV�+z <�1���g������=WIze�4�����߬��m��B���Rv�d�ʽ���+�*��ȥs�!UT�Z�[����[,,kn���DL�5�U�	��=�����G��o"��<'��m��|@��	�~�*��HW�_ix�� ��=2�9j��Q��wT���8�_
�pv�"
	�ɔ�>T�Wv��U��}�D�:y�u�1	V"��4.�N�+9Bt"������]4��?� ��k�~M���d{.s���&����``~;��s�p�E ��h<~��{UR'�c�1~2B����B��o���Ůvsm���Kp��n�Q\&�4V�Ѓ��~KCb8�B�%خ�I#4�/�d���f,�nϑ���XAP���Mɀ,ʌl��,��tLk���Nu+%W�����P�C��*q&�j�&L�Zi�ޗ���1 �+nt2|�����R���ѱ�2����֖�u���ԃ҃�h�^��Y-̤ ��xմ�t�tH��my�0������}/�Kn^e=�������^�g��:S5���9��䃟6���I�M.(\�FV���ڮ�+�vT��c�kб_�鐌d��5ݟʐ��2��-�
ٽЩ�����Q���<ƂT��:��}��P�pM�n�VɍT�7d�H��^YG��f�͌��B��Iq�ůgOT
�k4��C.����G��*?�ylP:���)e�8��r�0u�!"ӷ�N�[c���W�ftx�,PYV��H��C/Ƕ_�/�ʒ����܇e�\�CZ/�l�\�~[o��L�
.���QӚo/o����T��m�
�dI<`��AYܘw2�{|y��G�[5�DV�l�})NСm�V��>�t��M�t=D�.{G^�	:�P2�r$f�6��{j�*JTib Vii?���;|�d�ʇ��x�U���z�6&���/��㜽@+s�����kq�_��r������j�s߁.PR=����x����[�>9b�$��SSM��nm���QN�.��E��p" u���E}.S&�8{Yo6wj��e�{�S�3����8� s+\C=�XG��ܼ�Ll�!Z;ݷ� �dŭ��Q�X�m�A,�W��k`�╛�|��wQ�3��������]�=�od�_b�g�AD�$y�_�ך�V�G���p�;PNv�g���q8wP���l�˴b{�?��pT��C�:��I9��u�]V�p�[��w�7!l���r��%�	Ez2г�j�ߩm3/���(��&.�.JB��H��5O�a.֢�R�:�j��v��i���^�}�.�3��_w�[����0�6)�T��#�d�D��:��7߀�S����⥒����iR ��E�ۦW�16!�~F��&��pjW�l�CK��d��%+����dJJƏiSh��A#�7�A�kM��w�B�e# n��=�7����:E(8���#�;�0ō�J�+N[�ؒ�a.��l��[�梌�c�['�D�@��s��Ii�u�����̩�	G���P 9��A�5�kJ�����m�i�e-�~�i���Pe{1�7��!���~���1D	��K����g$j[���yO��G>�ID�������3��T�w��H|:��봺@���6�6��� �z�~9��a����=�{�W�Ѐf����t�Ф&̝~�	E=\H���dr2Ww|x��%'z阙�X��(��i?/JDI7��_ݓ}9���v�§�:Be6Y���ُ�%l�����z2ϡB7U�J�O��n,��b%h�u��/k������>V�Z���]�;�(U��,Oi�����]`A4MG�>0,� %��[6X!�oN�8��x�x����眺��6�87�`"��)9mt4k{�Y1Kpc��{�l+�f��O��EH�*)4�wֱ�(Z2!��S�f
�Y4Η�U��g?b��G��[�f}�R���{:��gXk ϴ]MC�N�j�d' !�T��E_M/�/k�ʅ��6�j��<�1��.Qz�s��ㆀ�ը�Z���7�p�O�lPE!��k`�$ه�=ּ9�y�G����s��c�)�n�U���{Ȁ7(�6�{1��~�6�O>%�:�(�ux_����K�=lǢؘ#0�Q�xCC5F+�tw���N?a�1Jt(@�Qޠ��`m�O��`���8������Ѳ�K{� ˸J�]{I�ߔ���tNj�{Qx
��d�i�S����d$Т�^5g�H��)mR3l ��k��IGwU�q�6{�PѼo_)�xڻ��N��Q����z��uC�L�Kq(��Eh�ʈ�$����gr����z�
��C�����ճ6��]�Za�|�G�LJ��|x.-��(�Ϛ���ϲ����pz ��Q{����TXGυ�?
AZ�,�A����i�T">�0��]a/�xz =�GG)C�V��4�.�S��;�Oտ�#���]��V�:���mͪ�� V̦y"���L�K?�<�������PjI1��4���=ɺ9��I	6�Ln�-����*�Hr�[4&�B�M2�R�ʶ�UD�B.Y��er������I���Ƽŧ[ϯ�t���lI��L�u������O=��.�M�a�2���`t��_h=���Z¯zo�&���[h��XG��	��|��g*Q!�plYު	+��{�Jƙ~?��/:c][#5��7��w񦺡��?`T��j�����$u&V�>c���2�+��r忕qF飞���'Qqbut�Q�LAҗ����W���p{:S_����]t�lP�Y��3�eI@I�g<�D������m�
���8h[�c���.�<���U"@���ҵHc�fX͹���j�"�k�F��یV�Հ��(?2��,~�x�`�����c�q�����p�G�X�{��ے�! lz�%�Ol����Hp<�ڃ�o�T��XfЪ��>����(���& ��E$��J�[!��Sal�lBOCqg_A
���j�1Q���I�3�[g� �Ŷ�{WN�=d@{��l�R�^���wN����h�1nV�M��;�w�;ܯR-pڔ� ��ے$D��C�������v����)U����9�鰭�`��ԉ��U�xI�5������D���f��������&1���Ц�,:��=~�	^Z���uʹ�P�=I�ܐ�S��U��&�\0s�',���Y}=�7=W\ � Y-+1��҄���v��|}@u?�'��j�@jt��}����Y�s脌�x���"B�AhΜ�2
��_�9�o�V�C(~� 6�dA�_��"��!kIQ���S�|�7[ST�H^���h3\G���}�żv?���&�6W�5-�Άx{�m)͖�ң�*��`$��E�"+c$x�i3"�ST�m߭�c �]��5"�e�<�-J9�ɴ�g��羅Y�z��3�u�l�a2��;��,�/��]1�W�|c�aa1x�d�QJ=	����h��7���œ�"~�Lo�rE~���{���;ڧ�"��*
>���uj�O*@��l�k� :tx\�M���6����H�ҙUKh��Әq�>7���K��yA��nK����W�1A�:te~�Q�˫F���]�Y�I��(�ԋw��� �_i�m]\��^��8D{U%�y���(���f/܌�H��U����F1�S��"Z�efl@}i�Ѫd5���9*�?��h�\�a��*V�68)�S�����B0s"(���N���}�Ⱥ�T��F1�d,�}�Wt��z'%�Q��9"#g@�̚�6��T���}6�r��4�9�!�Έ2a�E#½����1�뵌J4I|yY�`)=7��m�1��MAJ������ql�|
|����ҠFaC�0��nd��&��K�>Ɨ�.�j�Jr��V�Y�Yb����p�6��!�> 5���sK,���y�\���!C(�kFM��ł�U�����)4��ؠF;����8��x�S��8�5>��*ђ&+
��/�z�abK<�3���Y8�ɓd/�+��������˫YC��'s��pm� ��	i�b�?��?�\�K�8	�}��^����ԭ��%� ��A�.^{-��d�$�կX���}�jL����=�}�ʮ�O�/��Ç�0�8�ň�W�+�]_�����?��p���1E�o�0����Z�͊�^����H�n�Q�0�����dc'Ͻ4q����I3��(����7�<��5�v#ף w��57��)GQ����>�����^��B"���C �O$Ͼ*q�>f�����l��S[[�M�����B��̷�@����<�t�R��R*����Ņ�BP��Pe"�<�'e�>�{��]�e%�j�����~8����!��N�4Ŵ���&�2�m��^��&?�baOQ?Fg8�X���/_J���_����U'r�����H��ǩ_�"�@�� �"w#�0�Z���~%ny�M�[گ%���n�NP��J���hf1�V����v0˟G;�<(�-I���d�"�#D#C˪ÔpKoZ��\�f�Di�s]Y�I�k��c�A���2׸�#���������&�]e���CTn���x�7!��������!�.�C9�U���HL���9ʐT�(��p�6p�WǓ{�Koɉuc���Ӕ�x~)�{p{���Fp
�\jRe�e�c���t��J��NQE��{R��D����!���1���+L>��х�O��o�ٽY��>Y����1���X{H	��a^�#�q���r��p�+ݘ���Md�l\��pd�^��F�� 3��gL�f�_C��@qH�V1�)����{���bY<��F���G�o^ƓU"VM?�w7�F�O磚R'�={ާ�Lv�N|В�p�y�D}@���ʴX����C�b�$��41�o����R�g	��wሿ!{=-��(����)��;��$J8�T��
G^j�{�BU�.���P>�:��k��Py~I��w��2 �Xg��69FD��]�d�
Vm+�L��X�%qh���)_8x`O�1�LUڅ���i)���IO�X||��&���x�鿥ܥ��V�L3�����fal�'x��2j�|��`ǃ`<�^-ZR�����u�bZ$d�>m�����f��t��G4���� ����������ԓ���ϒo?�26-h.�r0�E���5��1բ�˧��d�:S}4٠\���/��A�����m���~tB������=��cŗ��|����e�,���pS=����Ӱ>���U���-e{Pj�6y�Ӌ��E^���s��f��/�+e����m�0Ʉ4�Ś��ۜ��C�ῼt�rч�9�d���g{ ���Y�.cb��	��d�m_{��w^b4؜r�YXl�%�άi�����|���M,F�}��\�K�
sK��U�ݢ3��Q�=J������_׻6���Q�?^m��a�i���&�n
�g9Wt֎��7��qԕN ������a3��� 3̢;b)h^�P6f'ci[���k_;��_���^���ݚS�^R�{��Q�F��BGx�1NBi�za
�>Ж���ڻ�ߕ��{"��t+�N���T�]�� �	*��>��b��,������}*����{�9�5p���W��| �7�=+ܴ	�l���8�*a��xݨѫX����,C��w�bH��*K����	�W��i�l�>��@���*/�̈�I?�������tk~<o����qH����afm��,���ϭ03��4&�z|ojC\�Y|�k���8)P����gq�@�	v$b2�"�%���>V��k��+�t��k{�Bቔ�uV�E������Ǵf�p(�1n�hhq���=@�����{����ɗ��e�/3����l�闣'j�O���K���m�~#�^D��+��4�n�?{�����_�J�]�3
2�9��i��a5C�&f��_�<�s
����%��h�	�c�=��0d�~�w�u�+h�"	�wȍ��>T�R�>���H���k�u�諨܈��d��U�}�Cvqm�iK��f��"a�Ke��IԳ�N@�t���v�������MpM�wP��t�1�t�d��t �p�~�L��V-
)����
(<��r��v�&3V��G�d�>"�BةR�Qa��-�]��w�Ꮖ�A������%L�Xb	�ƪ�U�҇�Eu^������6�H�2�0�lB�
)�p�����Ç{�0��3)��������[%��Fc�B:D�9U�ٔ6Á� TC�;����[��Mk�7m?%�L���Ěv}N6�.����f�e�0x���=ZyL݃�Y^杰m�c6ǥ B�h���pw]�m�3�[�S`u`�N��H�J�Os��W�M�u�ϣ�7ڕ=Xcs�]��9�>�tVK��oq�I��Mgߜ�g�@���fL�Lϫ�y��G��y�b��ͽ���TG&#,���e/������	��NK�Zc:|���-��k�~M��Z�u|ujR0�R�XZV�C�A����F
��ۺ�p���y/dQ�QT;2����7�S�P>�2'�#�ܒ�2�((���26Cu�.8�]�G��#mg�i�.�ؑ�����E��v� �#�����W-�j`��Zy����_�(�
�j��2ĭ��f��R�A-��J��/$l�����;p1�`A�=,,1�o	�&�{d��%�@�6�T�(�L|J����1<7u#�AT��A-��F������C'�s��,�~��'��ee�Bs>W��e�BG=�S6�=F[��3��H��9%�E7����+�4���<yr�~��	F�L�/@L�?���?�S	_o%�˝�NŸi�y���s��L0��������˘�f^��a�ёtlI�Xc@�I�~Vj�`� �U��Y��
¬Ώ؄�D��2-����i
3y�q�w����ɼAQ�����]߆C� -T���P ���e�'���b��Tp8�L��6��f���!��K��gl(�^0xrq�8��
W�c�W�KIv�w�����D�Px_u�q������>�_Zao�l���U�ȧ󇂰�p��VJo��p���`u�l�!s(z'`����=d�I7��LM�y�L+� ��(�������