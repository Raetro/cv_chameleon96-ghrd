��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0�����=�e�%�i~��Pt��	�)H���SR>��*�ptY�/$C(�Bl��J9���=5`����sJ�������y��f[7�]������2�K�C���T�wE��y>���_�-����O��Uc��׍:��2A�-�#O���x��m��rh4�k���y�'AsO���g�$5*l�-#?t_��������n9z��yAp@�i��J��Ô�.^��������{T`M���ǪG���CyֳΣ����ec���ʩa�Q0 W�q�2�$��{ٖ5��i�S`���b� 3�on�L=��YA|��,��*��s?y�� �vv�n_%����UQhj�7t�A�;55>�Y�%\�M�S��fX�zs$c�B�+�G���ɧ2���ۂ��:��@6��V㤻��z�C4U^7��vF�ց��l�\�/j^�5���:�JtHN���>��5*}�S���@_�['qH^�pLQ��/�e�L�����mW��n		;���H\(Rg��"U�9P�2��;���H��Ȳ�yXW�QD��t$����u�D� #��ֿׂ�����d�$��R��&��u`��F!m��Ų��s�
�Ȳ�ɼ
�V�uu,�����	<���L�����D�M>ܡ)�&���!2�O��o�����c�pٙO���Vq��W� �ꟻe
�u��f_D�H�Km�I�N��?Es5���R��נ�W���_4# �^�ڄ\?��!�{fy�BC����s�Z!�	B�!^ �w� �-C/�kH0w*���͵U��y��wP��q�������	x�3ˣ��w4���վr_�I�H�t�EO.ԭw��_#����-A�M�!K�n�t��_�0E?��`N�)٦~;���'����Sy��u�,�i�۪�,i(��/��$�l��J�RdR�63���w}L�؎vSK��^�p)��DΔ��=2� J����n(ow�TE�z\���O�}9h�SD��U�09.+��m���mtɖ�͛Ƈ��)�&C��� ���|��7d���V��\�K�P���!?N�r5
k�\5������,��������h� �K$�Kxx��xP��"&>Z�5��8@|i-�#]8�9tR`�
��}�̻�L�=���g|S��y:��u�qTN�0�{_Z<�o�o��j�����}8'�HO�n���l����1��o��L̳}��8�>e�����$��MR��TJ<����4�����b.YqI���H4C�8"X�5��)cH�o�;6�.;��`��ir����FYg8t�W�_��rQJ��������a��pc�!(�����A��\�H�ٷ����x��`�S�������ga��y��� �b��iy8�1�e��Wׅ6D{U���e$���k~�L�ѝ�n�xxoOI�pB"�c,S���� ;xg��t6+��'��
Mx�H7���⟽BF�:�ӌ����#��q�-?�*����W��p!DY6�Y�ZK!�Q��%QU��M�őg����쀯��A��`�a�L5�E�������k�	K���hy���ݤ���~���Y"��y(XJ��4�8z���4�^rZ�C���YN3˹��r9�1��:?���Au��@2�����gR��%'inC@�j�I��xz�]}Δ�d��k��֨3AtZ����n�ᓺ�l9�U�41�q�Wk�u<��G1?]o��d@j������B���~�V2��KpqJ��{]R��es;m/5:��n�)��鬕�2exUp�v}?�I��.�_)���C)c�FBo7	�(����C���=��Z��g�� �(��D�P]�z)�I�t+>�A����.�t)xq�3*!)f��L�n%�k�o�W������g��i��d�o���F�{N����QY/<��.s��B�-GZ=�i���k�%���G/�J�s�O����i{�A�!c#,e
���	���l�H�u���U�2S��5͍w����¾��D�}�9tH�~����Ýd�yi�D�&�d#�*��)��ًaphM��I������n��-{�B0'ѵ��85�D�&��2���v�&����ur�:����1P��O^��Uq������ib�>O~�E̌����f��������Zט��O�������;g/�y?p�Li:�lqƌiVʉ ����� ����8k�=��{���ع�H��
dO�ʞ�ւ����D ¡^H��,}��k+��;x�$��� �3�9�=pvi�����unv��7V���n��8���Z�S,���+���l͕�"�;��_3h����~�٘Db���j����gdrM*�j9\ֲ�7Pg�d���r4cl��c��G�ɣ��l�e��	�� x����|X{���0 4-
��`� aU(�%��3��Hv����W�jfe(����*��}O.����~˼�6��l�i��N�^���Szv��&�(���֗4��xu��2	_iIOC�G�y��a:;���-/���^V+��nQRۡ4r��S��$�f(G_��?c>%we����{�(ժc%b8�1���O?|��"V�c�`���{�Ttd(����V�ߏ��l��X�<x�!H=ߓWcx�yeUW|`?��Fn���&R�g���H��Rx�>�[�Lv�����o�0������g�CpT�.�����W;���d 	���`�0���G�A�M�:Yn�mT���֑'���H����� 6��{���.t�G&������ikNu���O��S�h���ĉ��_�C�m�����@��\̋9�̓ok���	�Q/\[&����m���W_����˹B�4�/�(A�%����<9�r���,Գ�*`�-���%�gHb��j��
���2���'?�����.|�~7��+CH6i}uj�K�Wn�4�8�ݷ�
��q�G��(�Z{T��c���y�a2/[JMݸ��n�^d6�s���YZ��s�_>L�@=���L�����Yd:y�k��zJ�N�4�Q��T�Gd�k����U���,�pp里UZ/���_�E1�F�n����zE��*��CI�pH���0��\\U�=5�q��:��wFX�?ݐÿfZ��ކ�|h}ڹ��v��O��{��˖)R��7�$����
���E�/<'\1ڍ��s��A�z��|�M�̋\�?�]��Y5�.v�J���,����T�z�7��:�)6ad�!q�O�V�vH�}�H��B��J��
���1�9ո��M=tD�T;$h�'7����S�'�
��vx�d�	�>�y�D���qÒ���#��?�%�.�Ϩ2?��C3rX�"���m���W�\tNa�[�F~(�#��֛��I��������WӸe�\����e��x2��0�M
�4�ל�S�����8������1���@hxm��gN�~+�p8]�݄��f�4`�k$�˕t:�V	6���Ϫ�
�X�8�"��1sW�W]֜�� ��+�^𗷤�!�wc�������$m�rMU�֋�b�poI�#��n����ZY���#l��(�Ϊ<-���M�M!8�W�B�69u(�3k�o�ձA(�Py����@.��Q�J�a���=�-�����u�J\�+�VB�����Z����ao�
7u2� �>pR�L&��R����SUy�aw����~ŤC���9i����$���p��Bz7Q�Ȕo{����@�~�����2��� G����h�M$�
�����5E��H|{1�ȿ�bM�0���~bq@ѿĊ�,�K��9_
��lH�I'����BԊjC4?ӌ�:��B>�5Ç|\�S('0O�3
����1!'�Y��(�����$��a�cu9����Y=+E2\�گ���o>6sw�����@�6N3G����e=��8��5�D���^g%�����u���>杌���T��l� (��lx�+3n�#~47+�����?��Ϸ��+�Fj�(�Q����d��u��yIi}��ǢUn��kIer�t�N_!�&�ۚ�o?�a���I`�}�l��IM�8��Yj�s�����C�R�=>��du���}E-3q-��G��]u+'bp�<�#���f��'ٖ�tv�vv�'��-�m<� a��Bb)��0��~��!�D�Nz) 7&�Q�IS��2�������8Ya��U�P���� O^ۮ-��4�͗�WD*v�Te���;���2� [���%OՊ��k4N�]LAO��Ef^�VVm��] Թ��I$z��f������lW�t$H��ǽ�@:�v�űA����{j��)���Wx>/N]�e�V �M{��Ym��B�O=���?I��jB2po�.�������� D����»��\]�M���_fֲe��;I�G�����/|C�F�ܑ�=k��e�k��z{7�wl�Ͷ�J���4�Ӓ58�e+P����t⃗f0����$�FRG�5�`�����h��ALJ��4��
1
�&�/�Z0ȉY��#wb ��-�g+��5���s�[z��	�����⟖��<{f�^��E��[2߫��1�>���W�`�oF;��<���+:�m��2�s%F��%�'섅��3"�M�aS�G�5��pI>��hxx�=��]���vf�=����wE@�#�̳Z�2��U����o���IO�r�	��,�{��9C���������@�g�����f����j��w�}XA����b�Y�3>6�('#ZE�T����!�^��[
]������f���9�-(/l�s�Uڅx^(�*�Q���;����A�:�(��6&��(�Rm�(,��t�wTn�oR�F�!3H�] �^��n-�ڄ\E�;��lD��?D�E���|]r�M�vM��>�P�K�7(����8Z&��]���\�K��0�i��eoW�L��	���#��)��l���Y���#FE���]��Xc�`,��	�+V�#F��۾<��Ƌ�ׄq���%�5H����˵��\�,i���D����.x����PH��w��E��0y8#�:���fش���Y��q�&Z~.�HC�������~2j<�'~qB��8D���5>B�8Z/A����M,3(!2LqCۆ��fV��������X@^�(���ml��mI&F[���m�Md�7���ޒ�һdq����J2#���6�;�7����w�`i��G�%Ew�p�� �<gh5��b�5���a�g�g���2�Qf7~���ϻpN�W���8��S�r�����j$L=��������� _��$]�,r���mHb��f��5/g���p���H��n�w��q�-Yq�W�w�G1�����1��M"�w1�_.�T�y% '
�Y���Y�0��.gG��[��,����������j���\�'zo�1	��ohzS�˸��x�ן ��� � S���@�-2�� v�h6Hv�(�
�r��t�$@{7�i��Ȣg����Y�ٹ��i" �N���'����#�c�=@S�N!�OU�Q8ր�|�@37�}�`���z�4Σ��_�#�=ӝu��b'{��D"�	�B�����v=�B�5�a'���f����ك�h�@���G3��W`S����fJ�n<�؇U;�����Q����XvYSvπ	�G����3\�k3������?ƕ������aD�j0����XT�"������rz����Cd�~��,���a�o�x+����H�n�J�7i�։62�3��bC2�D�5)%������)4�D�љz6ɻ�u�e�4��(�RF����ϵ��-P���f�#�&�I�����1�*��\溎ILlΥ�J4���i�����<�z���L�o͠D#�1��l��?O��p�*��p:��K��LRe:Y#��3�w_U��$k��F����M'��c�����I����y�v ��'i��rk�&p6(w DC��S���:�rr��2T���:4�(��&�H���V=*�%X+ a(=��"E����d�ਢ
:�8�犒%|��M'��Ѭ/mu��1�,d�����=�Cֺߐz�5�[8[�J�z�����8����6��h��a����Q�JH�`*�k�9���r�iK���ebpB�Qe ��54c��@�?��p2�K����%Ik�d�]O���Þ��ce,+;��"��kZ���{�����1���y�c��n�o�?S34+w,w<�lb{�0�F�8���:��^Ni�b�v�No���DW�*���o���Y��9���iGa����2���$�Bt��he3�n[�t%A痚���9��3.4xP��/=��S�&"�3G�g���Kl�Y5�u���e���8�pI�[$�j	.~S��H
�H�|{�H��Қ�s B��)�O�Xa�%���Ҝ��3�����6�-~�A������W׽Mo���*+Rö�/�/)G��s�b�[m }7���s4�&�	3nR����C�D�~��N9�6�f$�����3���j��������V��r�M)Et���}&�a�����d�?�.��B�W<{R]'�&�1��o y�N0e�f��,��dI�~p�Qӟ�t� �U�)�콬Tr���`��L��F�[�o.�� �^1ז��4�FȐ __��"�������oY6v	��[�R{��,�q$*C|�C��JVJ��1a:j%�V'k@������3���{wP=��):����j�=����0ʳ<��*�|�\�T]i�i)�j?.Ü����ʂ��\���`����5	��7�>Eę�7�ɍǒ��S���Mt�4h�9�ʙ#W�>�ڈ[���˛���)X�m_ȓ��^��.Ȣ�r��E"z��!�V��N�8Q���)X!��@&V��FJ��9���y�dX�E&�]Kw�'�#1��,>�֯�:}΅�	�c��j�!{�R@��J$#J^�H`��TP�	�)�Z9J�PXն}�og)���s�:dvO7
e�#C�b�9@���s��@�G'�A{�r��g ���'e>�Np�<�t��wW% �	�w�Ʋ�[���w�ޝԤ��-�ȋ-�"Z�*�oCu�rȨ_kc��۵�8�b,���7>���NtI���N��G���[M��	���j�o�?�ΔE�ΦӒB����K����E��b"�B�\��Sʐ[��ݩ�o���n�l-�+���?��=yc�Y�v���D�2�!� `U�AG��䑢�-��٘����*+C�i����=�km�hZU!n�}���J��
uf3�X��c�����6M��
�0pm?�UC�\�|2�8¨1���):�F0GXiH���J���z�V����P�.(Q8�E#w��4�����0��2���7m�0��h�,S[-�����\�jR}�8� �O��X��_�����T�J�܍3e�j�J��!X�I?���K؂|�`�Й-�(�y������ec��/���媅����T���Q�'� \��~�d[`��؛+�w�4*�Mɗ&����q������f�?&��TUn��.C�}r(*~qH�R�a����������������#Zm�x��ܡ�ҹ$sj�/�&�ۨ1L�.�,����G�w��Q����܁��xe�ii�Ê!���0���(�3����ɗ{���������>��
�֫�0}�1���㣌�
S˭ж����������@�)_�D�G�+��H+�;�n�k~�`���!3]`�ʾ��K3� @��qQy��[
M�
g>�S) ~���*���56�7N�Cbv]w��kys� ��*+�@�`"P'J���OD�س���'o���W>�c�U�jDz���{8_�}���(m�}�S�����j<\��XX��7�~��N�]�r�f�f�.m,���)-�+��z[��R���a\?7t �����03,�{&CO��
�I�:�A�k�o��tW�J�d���`X���q~9=	e�ԝ�i�Pw�]�h�90&��Qqi)��򜼛���y� �RG�=(2�*
�C$6��5��qr�oZA���V����` 8a���﯂#
lM[4��B��3ReD,J���6S��0��/fzc:R�^:LY_̒a���;,/"
004�̀�
�+k��~9m�ȃ	\6L���.+��k����^�~��K
%�D̚�S+��:��J�P��FjI/G䠺�S�}X���P�L�2e���-��"��&�S��	)�b�C�=9��W��ޟk��o���>b|;4s�Y-I��!�N+����!��T������O����F��cH�F����N�]�:��{ɘaZ�8Ms4�4 OOؽ�B��|h�������
&l �S�U��,D���jah������?+!��'Yt}l��_��@Qʭ�@����莽���cKLVטZ�6gݥW���/�����*��-�ߓ,E��8�^�\	�ѥ�H{X� ���<�ҍ�M_�e�2�S�#������@9_�<;���Ҙ�� �ghZp^�N{���ᔍ@<��A��e�{��GDk�(���@J�nZ���(
�s´��1I}F�4�E����c� x\�;���M�;���>Ҷ�l�i�O�|T<���,%9HD�oH7�-���ԙ*�-j}�S���?Yq��޿�.�mj��:`s΍>���뺑$j\�,�V�?��qj[�{({~�qL6���1S���C-=�SE/V�F�4��9�)�T�0m�>@�@!<�;'�
�cPTJ>�c�x�� "F&��������'�N�H�>B��wyۣ�
ro3�Ŏ�r��V�X#�����B�6�=���}&�X����U�6��ӌ��\BSd.y�Λ���U��dR0\ʵ{�Y��"R�Z7��Vhz3PCm6N^��%��SXV��tz�S��o���M@�Ģ�ݽ��ـ?ſT=�.�b�>�LL�'�J�����;1��p��=�I^~�ք���	����S��� ��h���v��o�V[�_�D���,<f�ڔ,T'���kk��o��r�P��we��)?c�A�7w�349���s1����t��٪l��4�FD5��M��LB���"H�����@�`�ƔL�_?��"��0���è�v�E�H"�p����o.���%�!�Kj�N9} _���������9��mc�6���⃎��,-��
�9ߺ{)r�(席H�A�����7���
����:ql��[���	 L����3��-	e�o�����ˣ ��T����f��mQYsՀH� ���T�5b����~ӿe�쯆��?l���5",b�9�a7�!�R��