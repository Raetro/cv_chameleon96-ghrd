��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��l�����f�J�éy7�=7?�w�e���˦��X��(|�EN��:D�*��{-� {���hEې�_�p�P�Fॹ(����ұq���[�A�

��я��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�s^W���0A��.�\����4M���ƥ�^|Q� oh�S��4�Id^UE�
R;WR��ΘA"�c��mK��w�C�c�L�s��8�(g�u�5j��nW��b����p���H�ZI�PxUN{���рAW�(6β�63^��>&o��h�+�	�UI(㮮���L���}�#x���y��o�-_��S��{�>u�*)S�^�0��h��v��C�}S�Ѯ�R-�ܬ�ji��$�s�m7��'?l��cPc���⨠�lb�Zָ���C\��Y0��ۺ�0�z:����Y_RNl�
8�.�5[���f�U'�E�q�;n3�T4�#��PҺ���=N�)
�<�I��������k�`���*�*�z���L
��F�.��F�j_�f��e�ܲ��Y��u�oޗ(w(}��X׶� ��ٿ�g��Yϕ�FQ�R��p��>���\%�O"� Y�G~}���G��p&z���e� "������M�_�Dl���~�͠=���]$��.��KVI�jM��D�U�L���I9��+gf#H�nA���ڿÃؕ�3,������l��ZPq�mH�E1Ʌ8.�iՊ�km
���D�7�ݙ����Q�?n��K~u�P��\�eM��mL�Wo�)o(B��*"��9�p�Js�9���B�'���x�a�(tɹ� G��<����x-�mn  �����wC�5���
�~=6	k�ts��H�H����@
��P�����-�u}���}��rv��B�^�cnMO�Hp|vY�p�)ߴ���i�x�+��!ޔ
n*>v�)!�����%�$H�_d��@��&�@�A�1K0�C���R!
DG��fř���v�~IV*BC� Lr�'�%�k��'�|Y~����6�](������~B0��7�N����z���oP�]�߆��!7���u�PWA�M�wl�n��jX���s��}�+�f�ӫ�8�L�0>����-�	g��3Vޖ"ȯ�`ƕ�f���y0�n�qU�b'�n_�����bΘ?Ti�L6�1�� ���9ݟg,z
8M�r>����VYK��"9�4�m�����W}�J�]�I�٧�mG_l�>S�8B���r�T$�����t9�[l&�.�����Jl l:["���{�q�T�$�|L�ir`ŊC�C��H��Gj7�pJ�,��A���5�f�[lf,�+Σ-��g���i���K��>X�l�1��Ņ�(QKV�_g�m)�8jO�a�03$��}�2�^Z2��p�p&$ej�����Rj��f��k��/�:OZ�u�MFY��F�f$���J��� �y#�Pw�B�S����F�B�o�hJ���aH�q�����#���,P��z�%[�hU�����S�b�I5n��t/�g"�	�@o�fr��c*�b��/"��0�U]�֠�aI!i�u�
��TQ�N'yb��g^���u�]��4�V4Vh��FoXy�����o+2�۪vkC�>U�s04W�c+m���ஓ�ܩ�[�	��<@姧��*q�ͫ��� �c�򟬃�4�}���*��gԏ���	�~^d�z�f�����U�++fs-@E��y��5H�q*�����j�}�̬��D��k�����֣�s睦����W�GF��<���i�axw��D���r����<_:�AoA� 3Oxt�q�G!�c�b��q�l����ś�'�����[�jk'%x�Op�DA5|]F�7e��J������
qAގ��1 �v�W5�^DY�UR��F���L<�>����eO�`�P������� 8�B�e�1�d�.H�/��GB�a)8җ+<uRy'&ړ��]{�=R����]N䧶g�2���%w���Ȅ��s��	��@z �M��y��q�\x� � �u��SN੔��Aۇ�ߥ}����m�0Q��Ь�C�v~Q�����l/8�,l�!r������f���,8ӝ�A-H3��h;�W�=�;��Тg|�_:����/ �yHFhF��=7��������c���8� �.K�D!��n4����nW��١�'��3/t��S:s �t����R*d�� d��3�}ý�a'�J�pM�Y�GP����ư0���ޫ�	?v���.�g�,*��r�kq�M��B���M���6������h��Z�B�r{�z�%?W��$[����;��{ԿaW�/h��՘nq���=VƗ��XV!�E�ԞM�_6M6_H�n�'�i�'�}����u�ӦK?&��31g����O�:D,��b_3�xŢ��m�J�r�߶3.����V����Js�����	:e��u�Cs�^x�l��9b_Q
I��pL��Ϲ�C��>�����'�,�D��B�ř���$Z��?	a%?�E~Ũ��*��9�o��V@)���l`h�x�ԤΩSBןblV*�U^-����p�͕,$Q���\
9�O��}��}NuT�"1�f#�B,i�������^�cF��������o& ȷ�Q���Nu�4i)XqPj�dI}��/�aweد�����؟��pp�x�B`UR�����Nx�T��C3Cb$�jۮ#ۑ��3Q��ll�+-:�?�o���^O�v�[Iݔ����s�A,����6Ot%��G�]pF��H.#�Vs�����|H��{�uF�F<7Ϸ�SfڳLV9_��.�E�j�	h
�!�h��M;�W���M	0̯���a�?��r�����2	�ԭ~M���H�X���w���7Z�}�%�W,&��1)u[e_n$��B�6~�sVl��>�����.���������9P�\:�����ׄ��p�f2�E:1��)���+v�Ҧ���ٞґ/�0r��i`�P7�Ũ�4X>DU�".��Dߢ�;�j��.Y���P@ 0��m��ɘ��Lr=;
���G{�0������HlV�G���Bqn
�""C�u�4���'�Q��ZD�H&�׻K�ͺ�G ҦO���[�q����ۿeE8�19�.�1^�R���#��V��p��-\�c��3�=�{��1F7�w�f5w�J,�������a�&�F��p{9�!���(<|�ws�8�wCĀy�����c3��&�s4�- c&�Xo{C���\M��rB#���@�d?=2�Lx���pp�@�Vk�3��J��<΁�Tvi+:�q&?U�{�]���]���ci#$L6���_Z�����T��ݲg�#��Q��8�Il5|�+���'���r*tCIE̞ku|�Sz���|_zm~0߹��i�Y�Ȅ�v�� p$�	Hܟ�s��q{AW1�RPܯ|H <|�D��Zb�~�U�^f��$̓�yX\�1�3�T�C����V{��K6�k;���OON�=��rl�Xq'o����Y�+�,���	ui@��G(1�d$����g/$hr�k�S��N��H��_�Cޚ���K�����"V\%0)h���Ok����Y/��}�Ŋ��,Ēt�6J�fY5��H3�o$'��f�F�% ��+����;"�� �Z�Ef�x��֊@Q���.L��,��6R����)�[�z�x&�u��pq��8.ew�Me.�J�*���ړ˩�:Tx'��@8uQ�#L������ȍ���@l��a��1� �d���st�m�x�#�d���3;�ȑY���b�~o`�� @�[�4Zϩ�I�� �_Z�DIQ7|e2}���s9�=FyZ�ܓ\F����0�?�SI�4�2cq�uו X��A@��B꘼fle�Kq�Q�L*��ِ����ߵJ��[���H��"�=�Yų��k�ȧ�/ik�~��};�-��.�zb�
�2N�Ē��Σ�؛Ӌ9����<2�������]z][���£-Mƨ�����p,á&�	�~8
��U���(+s���g4)m�8�DO� �d�
�y�Ԋjp�m�#��NՁ�:��K�C�H�2;F_3�-�3�	����\������r����(*"��&	��"�,e[B�j����f�pgT��O���ڜm��o����nslw���~���%���<3~��:�*�H�����Q����}$��T�W[��s��
�щU}���lR���XҴ��w��*N9�B�t� f����HH$&�6�����}���5,��D�w���ƣl�Or7���t�ƙZaш;���%����.�y9�����]��_��{�A!%�R���$|�4/*Y���]&)��6|�ǳ�&%�nΖUJ�����@:F�_�u�"Һf��KH�$���Y�͇h5��hP-b��"#֏p���)�FG�/ �ͥ��V�A`�Ÿ%@�li��OK�c)%e�x�#�9���>n�yo}̉��`�P>���=K���7��2�Gr$f'���_�5��60�G�����k7�����]���������N��D����d#��b._��$ ��GZ�`�d �E�r���K�Y	��f���*Q���A���r/�CY�M��)�:h��<̬R$Ju�V��~���Tz�<Ф&Ń����Lg�`~^y�&_�e2�(�C�1�\3�?~|�%�:6�A@��Ty��_e�p�@�^-���j�`�G����9�u�E/�����	�����`���r�V0�i�'5���B���,�����S��%�6�y�M�Q?�8l��5�ĹH�m��"�_
��}�K����u�`X��!��QkW!_N{��]� �%��_k��Ot '嚤�.�V�g�s��;j��Z0"UT��z�`{ �k�ε� F|.�k7��3��0���n��b��P��9*)4�9�W�����Q})�я5��$7�}���N�q\5XI�!��E*��J����U�&�Ҟ����e��f��2���e��=�\����%m���5�aO�!/wy���i�ޏܟ�0�=0��0����f�|����#����'������9�m����} ���<~�O�C��U]�bc��2 8=x�P�Wr�
tu~C������$��|T�;&w�KL14�FK�ߧ�h�� �3M��&���q�'@ҟ[,?<{���u����I�l$aɟX��E�Z�K�
[�d�&�����g�C���a��$/X�n3���z�
_*Fh�=r2��UŢ8�A(h��#�?'m��ܢ<=�:3
���|`"ĕ���Gs����P��}�i�����ަ�jcZ���%�������
�/_�L�ka�*6�1ګ�����~�CNc�o�u�m��ca܇VĮ�B �󕸺��Cy0��F��C��c8�������0N���խ�c^����ޏ퐸�ixB_��������3W�τ�Q�12�q�%Qhp|�Q��Iį39�?Jgi����X�|�쵔?���q��I֑	pɟ1<�srf!	)�N8;�������%� ��җ�>JE�#������_��;�(���B��$x��<K� �fm�S�A#[`��MjZ���Mt!��@�
2LÈ�G[�`���D����x\��s�zF���5X�% +���σ���\������f_�{�{��x��υB�9w����S��e�!�[�,����h���
�Y��-̽t ���F��- �sƗ���X��J+(4����M^�f*����!�Q8Z!_,��e2� �Q'��������!>��u���X�b���^���T���~�ÅҐ_�}�,�+�yݑ�ʫ���K�ǇߝhB�?��>&>P�]�Zڜ,�u�{�M��.Q��8`FT�]�8-*��H9H�D"'��j	�2����P��ʠ�r�����ݭg��_+4�R��2�N�AK��i�&����ȩ���.�434�p�^V�3�E�����1�e?'��D|u�M�kS�� 5��g�F��D���K]�H��ŷ���R;�14J�o!'YE�+}��P�#�BQ�&�i����G�VH�ƙm�����;.9�Ε߆�w�oTxp4Sc����]y÷�	//��	B�pw��� 	Rͭ�� �=o�/6"�����*wQ�g����r���+�JT��W�����s�L���tAy�*}4��!�n�(���L�U�Z��1��ΨRZ��F��T���ƍ��Pk���/U�x�7��B��u������W���A��^�^.�d��YA���y��ሴ#H��-�?�g��)��"�L��&u2������,��v����Y�����&\{�S<�,R�WL��}+�Q�hD,
��i�E��9 �ey?���7��G�n���{ыO�jO�,����d�8g8�]d��1c�/,8}C^���A�{,9'+k�pQ/�hA�q"֪?D� /Vw�B�*N���0� Q�׶�j��i�SQ79����LW��.�Oc:�90$�X�EXtk���z	q���HZ��^���rMu�.o����~;≳_}�%��
�.� vnmȞ�N�	��P{�^�o��WWbnC�����8=��ؠTu�P�I��Q���Tz����OdWj��i%G��xH�j�9�7�o�"UG����6#��s�Nv��×<H
���3	�L��	�� 7�7y�6k��@��%G���a<��b妰ß	��V�=�)P�j�m߯��[�W5���i��%�l�+�2��gVy�`���p,�X����O�%��%�J;�0.f����A$sZ�ڿ�u���a^��k�gU?Ҷ�?I���\��Kn��[D�*�	�EZ���Z��2�����j�n�[�1:(nr󯏗'`��#�n�G"'���Xd㹣Տ?_,t������ӌ���4����c����*<-�U{�p�]g��kUf�Ng)����;�T�V�܂(�64�M�I�q���C�|=�ҳ�x��%n�6c:�;drb����q�FMBsWl�eF��Ż(x�4:�e��30Q�R��A��j{���?2�R�r¦)*���}�>�e��k�{ꎊ�c|��yXr}��os&�8�?�Os�ki�}�I���{�B�
���F�))���5Գ��(G�����4T����&Ls��80�0ywPrv>-^��@>�uJ��Cy���ݶ����c�X���8.<nT�=]H;H[8�)�D��㷥����5��I���q��K'%õ��N�@	n�y�\聓�!N��ď���jHmQ��F@�Y�^��IGE����q�:�ϸ�Vlt���u��@tI(���<n�d(�7�p���6M�skఝ-�J��Ϻ�$<����#�Z����*�տ�Π(!���6�s\�蔻������yEw���|�����c��7�Y'x�QLe/�yK���<��b��&�:� X{zԵ~~j\�	ZI�u�[���"0'J2>Ǥc���3����?�mS��	=��I��M�4Мt���[Q(u~'=��Ii/�@Cv�5GTڳ�V)M�/��ז�d���Ab{������G����5{��[yx���1m�b+�Bw���>�
�^�!NL��-�0ݛ"�t��:�u��q�� ���ͧ��c��e���NX���'7^���b��Y���h���m���b#�k���ެ�La�1�Ŭ, ɤ���R]V��z��3v)�(ܷMI�a|B����b�L�+��!�����߭�y�f���x��h�[A���$\��#�X���g�|�3�|�HXJ�P9��{�����[�}+
*�O��8)8���%�T��DݭmQ�v�zO-�*��Chfb�5���
."{��eS�1��r3��b��T��ʣP��"yT0�@dF�ֻ�0;��������p�Z�"p���b�Z0�_*b�d�T̉(L��Eϟ�c��o���ѳ2~�����DLOW<�PWp.���M][��yiM^L]�p�"��s�5�|�h
*����y�p�L,i1��Y�z���c�)?h?�����'�K��?�G����4�<m�W�z6��)OҺ$����un�|��I�>?ݞ<�tu�m*	@����5BR�L�O�+������=��/ZsO�W��w����KP��	f�8V�%ɋ��^jS�[Q�_�QS��Ͷ'�tɷ폟�<6�Q=Z�RP3�5
�qx��Q�1�x�!ďEr��U~��m����\t��f���
��c��N�Z�-?,��k�M�^O�����nI��E�&c_��o�F�~y��E{��3���O�^yǛ�Ǉ�gk���:Bat#7	����8����9!Gsb���"�p��x��-����|�k�{&���$�7L}�Y����&-���ؕV�Ai��#�l�e�I����,|<��j��
�ܜ�	>�y�ۜ�2hP��&M��&�e��f�<�#h��r����w꩓��?GxǄ�e������\��Ŵ,�D��;@W���Ւ���k����e4�l�a�	| fRJ}�$�DH��>=_��n&*L1&���ՌN�WS�\)�ǡ�ؕ��s��#���w����нx�#�@�Yt�90������,�k���=���ǔG7�����uM;� �|�p+�:�Fd Ӹp��7��mN?��_�]��xߟ���|kB[K*��$j��.x��ҥ�� >Вƣ��T�����pF�� � �ly�H�&>1�o	^��m�$ဘ	��Ml9��%��l"
3D��2V����-� 9�4ۿ�!e�a4�:���--8�p�rF��o% D�H��C�|�ܨ���O5���K��e�F��E:����j���D}���[�f|F���&FasrӜ��Bj�<�h:�?����J�ž[7�h��1^����n�@�
�e�^<)V"�v=�D�9G�U8� ��M�{u���=A���~ぐ�{�V�F
���VG�'���d����ã�ǁ�d��|S���;�)�Zgl����i���Y�J�N���E.�p��#!�Zy�2����.�2����-q��k]=�R�J�﬽I�C��_]��
}�&��BC�Xd�د�=#;c�����\[�����J\}ʿ,��<pe�pיA��p+$<�w�l��نjWX|�ذ�y��Xo��� dšť��1�Fx�xU�em�$��0D��xNdu��_��������pB�����zx���r�`�t oq��t��mI����\W��E`),G4E0�c� �C? i�x��M=��.�n��.����I1�^6D�Wٷk�KXcU�gwoヤ���S���02k��n��e<Z1z�����\J�� �͐c�R�;��bd�gl\��nE�l)0_ƞ=N?޳Θ&�@%#����Y1g���%E����2z+��:to�k�x/n��\v�Yd���CUY�lB̘�y�����'��R�nd�\�R�j�C�2P�VH�����_�,v�?��[ޓ��d4um4!�E��\V����c?Q�G.���#��\D+��7�dE�}P+JM[��4j����@��{Vq�J��ܓ�;_T�:�G7��X��K��&��BT����������N5�@ٰk$(���HV��T������h#@�Ӄ�1�PF��QB�pТ[�jA�8*��&�QfN�90	�f��{_M$��7F�3�Ē/��OE'��4JVKf�ݒ�ܫ4�E�
�m���r�P��U�F���N.��Y�m�.|%�ht?)��w������݆]��l��0˃~?�����g��� �2����S� �c�4=Y��G.>!���0F�>Yb��m+�U�Z�,�6���_|���|�S��s�*�(=	�N{�o��r�R���Jb(X,��;�ً�UO�+D�.ŸrP�h㞼?���M�.��S:�v��M%��W��2u	� X�"�B|�����ZNC��E���f�!�zàI$i�q�22��w�8� Fc�F ,]r�Iӂ��c�y�a6&��hl��@�x\S���i�����L0��նS�����,\�=��c"�^��Q�KO��}�&#x8�5�Piw���C<��G�9u���Ɗ�x�3�����F�r�7sB�s\D/�$��;i�i�?�i�^��V�5����x�
�Kw(��Dd�q��'������jhdt�%r������\��X~�%�M9tu�C����\�l��e���ڦ�	�	�{�N���#��K4�R}�3��lۭ8���EQ���#0�{�܌J��^ �;_cۄ~H��]�s�-LD�!��|?�
�E�=$چ���9V�J��<`F0��o�G�i]�`}���0��M�c�
��n�\8\x=��>m��?k�u