��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��l�����f�J�éy7�=7?�w�e���˦��X��(|�EN��:D�*��{-� {���hEې�_�p�P�Fॹ(����ұq���[�A�

��я��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���3N^eL@(>5큁}��YD5�s�v�%w�iڈ���5v4�����aԠ�b
��+e8��ڇ�!���#=X3S7�6]��n���f��q�fB/�RM���+� Q߈jN�������S�}�.x��(��hr+��x[1�k� �,$ʒ��(��������C�L�(�?V���nr��?&�?��|�ƪsO�x�[0/��.UN��ʆ�g���nE���"���ﰋ߽��c��+1A�H�i�502�)g[/�e�.ݰ�Z�)*����T�3�ie�()U
_\p Ⲷ��<1o��6�ٗ"�i~9��x�AF�3	4��4_P�s/��w�C�`n� uu�a�$4ڭ8	E�	C_�G���6�I����I�]�4�[G������C�+X�=�o��]��E���*كP��dS�'�(�^i���'���X�T$#;�M��K�zibs�bkgAXc���(�$%H��<`�|�{)�r4�N=^.��y�}�P;<�B���m	2���y@e�`'@��ѥBR� �@h�j�q	"$�vΑ>�[# c�3M93^*]���v⒭��_R�n*���g)8�g*���}��Kq#��d��C�jM�'p:ل?Ͽ�ǵ��__6\{��v�N}�!�EO�����oll�_Ǟa�y ��@�^0v�O���*�r�0��8�^������Y�Y��q��ZWx@@����4?��] ���`�n4�~M�C�<�1�F��E���t�:~��L纊���4�� p�-�Zň�%}�Z�Ӛ$��j�T2Z�o!�D�6l~Q��♦�$��2�$���Ľ���k@�K ���0d�=ZKI,r�.����!���1Ĭ~V�/�.C�W�6�6c*����3��q+(�������%OQ	���s�����^�d����S̾l�J[�q���sR���� x�Tx�GM'� *���"�ē
H�&K�,L--n��M�̞q��	g9s}�7�tG�:�G���K?a�RF�k �-��[�u��,dR�y��Rd��@8��c���N&$������q�4Z���$�sL��o�@�t��/B�p)�D�uio��9C�߆m�7����2^�{����$xn����+|uj���/��\����h2M��<8�lϽޟ��ߊs]w�w7��@^y�u�,d�Դ0Jxq���dۗ�[�ᄋe>+B�����!9�	~�O�H��M�3G��Nw%�]�hF������b!�8��p�נG�-��!E���x��yi�R͋~W�*�SƳ���鬒]���4,][����g�r�y#Lt"�������g���l/���)L?p���Y���5�Β#�5�p=�Z�c�t�F��qNSK6���N�6�N���D�S uZ�]"R����5:���=GH����g ���#W>�\v'/1����"������m��6�	�)��Q��u���FQ�1,ύ��9�F�* ��`W2F}{qԙW�3��� �Z�_�6i%N"�b��*�`V�����oy�a��k4�l�m�rO|%�z[iJ^��M1��sE��+���m������5#
�ZD%��
o��P_t���0�9j���I�����1�b�������ꗠ�$i�Q���n�"��!��22`'\���+�t�K�ؕ��w���)��՞rW.�%r�O������
~������[������BB�m�s�c{����TX�t��v�3L��c,]�`�?���0J.�5��T:���8�5��R�E����%`(}���^�A��#���,e�;��n�C��n	 a�@�����|��>;����Ƙ[YU9�1����3T@}[�*�U���6��T���^�����������XMK�ϵfD�P�!wg|�m�r�X{W]��聱)���3�ӧ�E�\l/TWl�,C,���/��e��3�B�n��bFz^3���i�߭q ���	9G��ē�0o4F���W�}�� ����m��r�@W!�?����;=]S���:a+r���W��a�͓��|��Kg?���#�\~�򬟌�:i
A4j��Ԛ3������5m�̝�Q����]���pCG��I2��2K��ݔ���],(!k�%���"L+���cA>eEDj��"���@1C�X��g|
�fG�B���ѫ�	u�L ((��2��U�6��q�d^�t��B�wܠ�#]Zd���B��/,����'�Q�o�)���ZP$N������R�+(ot��&�BZ(h�ʨ��iȧ�z�Ý(�o�}�4�:��l�瞧j�U����>��+��Q'{�K�� �9���K�og���`p��)����u�}�Q�6�v�孫o�#���T�%Q�tྍ�A9��3tNs��$�g��5��&1�l	L�<��2���Na���:�N�ս33�� 6ik�W��-��1S%��F�4(��I\��G�$��%�r�-0dEN�گA,�L�$�bYB{�Ll<�b*��,^.Um��.��@hA��YӕW�	Ҽ�~4��DQ���I�cK�����?o�� �v���T��zq�b�:���7b8P���4 ��61M��h^dyk�KMg+}'�Qx�
�=^A�u���^׮R���l#��2�wd�*֡v�OVD
ǈe��zר�`��h0����&���p����O�*�}pl	L>٩�"=EI@�Gw?���W���@�s2�e���r���p�bVڠ�	��Z��O;^#�_�4s+���6ܵv�q�8��Cg[�^y�k�E��|�ֳ�����HZ���0y�R�;��7���dT�?��ۭ��/��-/�bӸq�����	��G㏚��P����DP՝��ɺ�
�7�\B�EZ���J2�9&lf�V!�'��&�z\���8�]�Eȇl���d��53��:�^��7�.�9"����K�+OeN���PJ�����*�E����C�lpC�r��H�������eH��Ӵd�F���sg��i�Ni\{[3�u�-4끿��M�r���qA�\�
lu�,˂I	O��?k�R�+LNЖh�G��?b�p$����WF3,}�X���t��s���e���d���,ڡ��2 ��m��l-x�Į��v��J*Ƨ�d�eb��|^|G��duJc΂�h[�]-8��\<3�i��l���pZ��ӄ����E?�Ԫ�(��u��#�P���Q���L��VL�7e�S����4|M��O ��c8"��~ERV8��%'�1m7v^�gICӞȰE�&���ڣB�<�r=�H]�ҲN�Sd�߮ZL&#u����/eI��R!I���%ʵ���-�����Ҟ�Gp�r[��h�ZP��#P��o�9o�f�곭��I�ѻk��a[]@��k.I�Y	�~d�����#V�m���I~G�����l KǼ����Z#
y�R-9�/l/u=FF<w#����N���c���R�Sy���V�%O�^���,���bHC�:�����	}�U�.�?F�ݼ?��a<���Y��c �/!Xaڪ%F^�"J���5�Pr�2�RCc	A����M�8�=|�� &�^;�*��"o�kg��3ў�T��h�Bl]{��Ӥ�o���6hX߼� �ʻ%�
��F�|%U��"�O���h"���L��M���ju��m��!+�����Y�D�Y�ɓo]@ɡȰ��=̍��]Y/�O��
*��Ƃ3M�ԛx�F��i;؄7s>Hjh��j���X��Qk��C���A|7R�W���O��(,`����(X���/ѬfB7%�A
�_*= /��6!9�����]RT$@�̬^��G���V����U��o�N�Am-���E�@����p�ѐ�����!���E�u�E8�~Mw�s��6w��:�]5@�q���v�1(�#.�x8��w+�dk�5I�����U*�WC��o�;�Y�G9z�h5z�#h��E�.���Pu�,�&(��]ǡ������"V�JO^�C�L�l37z��D+�^��ۿA�ʘ/��ƍ5�z����d�v&�ڡ�9~8UZ��=��'ld���N���u�@��	<=�*I_p�������wu>nGQp\*�¦�Ic��Y�����8�i�\8�EO���D�����G�jU��T�������-�Q�d�ځ*�|������Y(�D8G�`.^
�fU�Lgڅ@�5� X���m�C��QP�-y�&}��\Jj��ogs�=Uy���:	:Z���mZc�'~*s,A���a�0�}I�����y/� ���_Nƾ��d���3C,U��{�����jM�ŧwu�;2);�t��P���k����]�la�����_��s�
� �>(]ok�S!���#X#���s�!?�B��v�-�pl�����N�? sm�S��]0,"ou�(?c����;L���J��5���!!G��hl�s���F~[�Xp���bi��tX[2�9^f�T���$uy���Î�3
�NMj~s�uΦ�|Ls��O��f�I@��q}�&b���J���CP��'��&ʤw<ҘK������p,;�mBe\"6ö̳��؉�3�j��ZS��q���`��?��D��ݑ+�~]V�|��J�6 �@�_Õ U$Ti���h��t�1>�x>Z�v�I��p煔a � ��X����AA��/5�c�E�u`d�J��Ԯ�hns��;*e�ռz�lqN��`���A�qHꍼ�)㥗C;�!5��Q^�v���-`�B�W�^t��a�R���>�+*�k�:}qo�ݵ	P_���"����6�Y����Ԩ܃s�T>��t'n�u�k�����ߚa��I�_���V�Ƕ�E����Th%C���M6�Ɵ0�3�"?���V$\)۷�O�7a����l[ą�g�:GM{��s�qA�\�͠��=<B�{ԕ$>'`�y��P`����k�N�oe��W�	_�m�c�2CE�*�%k����a�(����_h8�14��z8q'���
eG�����P#t�{���UM	�a��h9Z�C���}�jo�7���XYx��.UUH�-�ٔu2Ҿ=��q�� �>�15�<Z���?��zxC۵钚����7�\Y��9��z�,��1�}M��wʥ��J��� �X�}�^F " 5�j���?O�}^�? I��i���L+x{�	H�9q�ܟe朱���!~�3o�ǚ��b4��='��n���~'�{��h�!6��I�1� a�ҋ@<<ޫ�����sr/�q�~�5��d�"\%�q�4��:ŵR~Q�� �ѝ�,��Qy!0������W�̳�M7��=�sj:�85̫�2Z��.���>
5_*Ɓ�sew��Ke��v��s�zmN�!�ģ�d��&��i�E��&n{���!ƌ�v�s��[�%i�
�ƅZl1!��"�XteG��Ӑ����y X���=wA��OD�z�>�0!O��"pzb�-C�6��*>�)*2Xs�P�?�t;�>KT{�)Sd�&���x9=��i��s����,d���VEl��1���#x���A��[~�W��;�pv<�G����P��c���N��A���o�k�"c�)��s$X�Ջ�>s��xx�
�e$�{�{;�W�ؗ�%�x�H��5ͺ_�RGĝ�띺8��j���k�5�P{{g���}V�)��>��������ebKK�tx0F@b�|�c1:PΏ[��8���TK�6Ve�����iX��9>��I���6�M��m��P6
R��l����q$o���j}"��Hz���ÿeؙB5Ǜg��.$g#%4�!3��g��$D�1 68���r�	d�!��Ȫ4c��H�Z����6<�{A�:5�S4PN�[��HJ�|��A7�"E��:Ya?�(�Q��ҿ0m�"�x#օ�=f�r�{��y��Ӟv���V��p��`���~I�A��f�����<p�o��KE���:�
��c4u�����>�x��c��u�\�τG���䣡�?/�O���V1F$R�Qx~����"y�^�xIgo��Ϸ�e�!����>[-ئ+�̌�KB+}po���֦i���PW5C��J���ɟU�ZQ�F���
��U����}ʧ*�R�͖��Q�'A��.P0XW��mT;Y�~�O�M9N{*`^���܁�탘�d����}郡,�:�#�%�o�)�Xؓ�aql��굻�y�7�|�1�7��"�NF���f���Y8^�p	9��1��4	���D~t/�e�b/Dn����eƭ�t��#ɳ�IRY�e�_+��i��oo;g!2�ܬ�hT^��k�S��g��O�N���̸�&S�ʇ��9K�ͧ)��m��٘�t��a���4�wY��R���3�,���S�E�`&���L;�G&)��?��_S� ��� �Q���� ?�l�eb<��|	�6QqH�@��i&�z6���\���	'�ż,j+K���/���]&6���[��{x�8N�H�'�q�6��;f� �	@�k�s�R��-;� ���Dtױ|���*OA�j�������c�Ѐ)|:��"f�����}2[�1�g������)�`_6To7�v��;���Ma$��C�����6�%���S^j��z�%�Y�^�AQ��e�C�lA�H�ө��b=��!*�^sűNE1�<{�EJ<��j�Lڗ����d�Q�y�8����|-�����8p���X>�B�A���O��O�Y"I���%��>�p׼�Z��L�\#7�:kS�-P�_Brs9
��"��DP�=����L�kS����o茐-xW��ƥQ�I|�}9ħ�,Q�+�hP����b����H'��a$:M�þ/��h�>Yi�.�v�����Z�H��x�qw$D�
TԿʐVr?��,R�v5~�1��<����szXD�4�x���"���'�����ݺ5�R@��nd��;`�4J���_��i�YU��Tk���.+��F�?&�KE
���A�R��E�+C^��lr�%�RJ�в�ET�@b����+uz�f!�*VE��sZ��1����*�I�>&��	<��	���Pa�f�xf��@Oj$^�L+��I�Y��A/�c�1��M�5$˰jT�g��z�~XŮ�u�o�#+%=�=����ޥ����f����?�]�|D����SR��t����;:'e�I��#���u��.y�1Z�H[��^�d3st���qo������KZ��b��U�K㉏<��#�\Z��Ox_�v��~���[�9n�4�����c����V��חk�����0��i��YhD���Z�?�p���O��\�0B�M�ͣ��r��qM�Ap��N�2�nV,v��k���PՃ���~	���a�=\�ꑲ��X��<��<�<�}�h�jKIO3Ae�i__�|�`�v��
@�d��^`!��RF.�\�L!W�����R� �@������O�mB����>�3}K�����pN���!����Q������!xG��6�$dql"��A�����|���l�&.�+B�jN��[8�&�0���5<[��	٨�����lN�-�c`xA���YID:��#�ձ'k{9AXu��s�Bn��6��j��l����� WzT���N��ڪ��,B����_D�8��-| R�jb<�tO�U!��I��@Dw�Fݫ����\��?��#i��@4-��\n�\ři�s[@Vp��Ga��#>�������tO�aߏ83dR�BK��L�8_
�S��"�2����ƛ�M*h�����;f�ЯyY�cs�[&�M?"�$R!�Ί}_���A���n]��R(���L��6w��yYc�R��I�Z x�[��W���ZQ���"q��1z�}�I��5��},hN�{zCU��E�RU������\�#D愎~��N���i���-dv��V}L�$���K%�7����fJ�s��A���& �V3A+� ��)�×XƜ���8��S���`��l���`%gɬ�e֗J�ko{c-������T�lA��ӌ�]\f�J`H��!+"C9�ZuOsȳ?�i;�9�ڬ�=�[&ԕ䘎Чs�{mk���/6	<�����=�1��VC�ET�T�%��������L�h�?��?�QDC�=o�R@��I�ը�.���.�����K��]�,E�"K��ʥ��o�k��|5�V��F�ؚAU��N�.��^�GI���F
I��Ghh�������U�IM^3����ׁ�"L	��o����h�8�8O*:�ǩ@��N��h��P��`�d�`KZ+� @����/�m��c@>8k6v��S2,K��A�'M˲���v����Sх. ��.􈿡�`��+���:�)cQ���BH]��ĵmc,mGH"���7�L�O�(�m�'[�-\��;BM���L���k*6�	���[<J�Vn4P�f+�9+��@�$��C�W��I{�~  ��ݡ\�8"�K�NB���}��䣏�-⧘��s�hWM�ݢ�i4��F�Qr�,�gH��H=Sy��\�Q�����F5)m{r��Յ/�/$�k����C�ִ5��S��76���>s�08Y	��'.����X��(�i�0x�T�P7/����@(�c�_�&q�@��=�J�:<�"�Nд�^��L+�l����T�a�qW_���Dk#Q�/y��.�~LO��Ⱦ�Y&0��e8@7� ��Rӑ�>B���ek�¨�<�4%����A^5��qi��rxP�A��PW��TK��V�K
��W>E"Yy��T��&�tx���v*�&�f�A�Q�eL}(/q@H4Sw���ۺ��Eǒ�����Q��~L���#���q,���wGzlI��9�Po � ��Z=Y/��nC�>c�j҆x9�0���E1C������'F�W���w+%�e�G�2à�6D�0m�$p[�lc鵠1Ա������jr|�R����U�5�>����*�j=ќt0ی�:&�%��}�1l�݅o0�UR�:�er�|!d��(���j�B H��T��~ɼd��xDEV�&1�n�'���~��,�V��Em���g�k����{�iz�޾�!"p��E�p�q�{�AG�SE[�H&�*���q���"�P�m,�l)L�=�m��^�D��$2@>æ�0��Q�����ֱ)zV���c�
�����T]}������j�uK	�p�����bsC^�F0��:��p��G��5Lv��o�m3�,R����c���5��%*!�����>]`YT�%&SSa�[�4�vY�0���4<a���~:����{�]V�|-��B�����t�o�%�so�3CIS�掱�b����
��*mα�eY��
m����O�oQ�;�_�iq:}S�Т�!�׭:㰎��n��>�C�]��B��P1�����*+=��ͭ[�v/��p+�Cg�c]k1����>�yS�5#@��� �騺z��� �Lx�1�?Nd�>�y�rޖ`@����֦�W�R<�M!��֒f\�Xab��y� �j�\����p��uQU���KE8��H�e�3+��CM��M�C�|��_��j�>�C�6�?-�1̃���!ъLQc�e�&}��%�+���e��ia#ʥ�M��Q�ư����?�#��Ii��zE	EC ���1CK4 ��GN���>��1q�u�U�z@��vW;���}�2�Q�	$���ǜ�RP��0�YP`sB���!�k����@T.���k�3��5�o���m藉����^�㸵)�k����J��-�I?���W�^�l�۫RMD
�3��N��P
Ϝ��a�rb!a�������m���2��yE�w]w�i�@,>9\q���z��N�!^C�o�q��t룊ٽ"z*\e��K�335�tY�L��'nH���u�V<s��x��X�_y�1:�a���^Y�|(����CԂ%�d�O�r��4(刔(>#���ޤ�L8��b��!��\�*E���(��
]�Y��B���p�����ts3�J�x/8A�UF	�b%�_�w[y��m�	�"��{Ј6�B��:�Ԝ��(DN��:0��tx�x���`;���#� H��߆ �dm��uv%\(c��]/e�� 5Վ�?whPq��^�Hd�t�Y�/$��y��1�;ڢ0�N�%�n�\hT!��R�c��8���ՏvۄjS+\��U�qD����h5X�{��i'E��_�k|=��1)�
�]nĒ	�#�O7ҭ�N�M��kqjZ?5g`�B�����T�ʃ�K�=ڪ�'?���-�񀕚
�� \��1����Y�
w���)�*!�_�7�C���>�`�0��6]�l\|-Qo�/+�gS�jG��nNV��r׌���gҹ%5d���YF/\�1�f�^�[dYl#-���b~����!���-�̈́�		��(�����x6l�2����3].���em�曐BH��~��n5k�ަ��pƱ5��W��i��Ps��I�wp���@�����y�2�>N�o ip+�fs1���Ǆ�Jيu��l��O-{ȇ���<"�oa��Mkm��?�)�\E	V67},6 @�����gV�t�k�kc�5/�6{ٺ^�H�(�p+$�#I�3�R��k$|�HR4�7��-�;.�/��'��xP���y�z��go�h��j��N��2Ae{���T������rZ�#�t�A(:��-x"t�W<a�`��V Uv)����0�6�V��X0��,�8��I�o2'[�v�ծu��=`�RSR6_��yHu�����o�B���ݒn���ڈ��0}	�g9}C��$�%JKt�mI������,�� b�xhX�A�W�s[�A���d����1��?��H�DK1�}�"!8�4�򮰊�] c�3Y�m�D�I�2�C+=o�~f�qډcC��&�y`Z_��x�E��t�S��&�&6����b�W4I�yf�4�w����,7��6�� ?mN�qY���J��"Cl��a�9^�A�'űܘ�Ԅ!�ԗ��m����`+eQ����2�rk%�h�}��?
�TX@�l���8~.�*1��"�p>���L' ���&�����Nf�g�نy<��\��^{TDG��1�ݓg�����㍌�_��ϯ��kj�P��}"�6C��������ҳ-|��e�L,d�ο�.[��"�f��I�G6SP"�.5ӓ�}��	����f���!Ȃ�p��''EJy���
�����(/fgX"lE��8��]EPGq�y��o�1���?�u��H��e�>��l7êv^Ո�J��L����-M��k�@��"��S�� �����é��\��P��d�ZE !냦����,Γ^�o��܁�&��=��]�����:KX�	��ށZ�!���q7�GZ�ʷ9"TX��r9�S�<�R���'�Yc��Ɔ{l�<�~���{��.��<�ʖ�KaxC�j����}�R�ː�x�ҳ<�Ǝ�㩬;	��˱����a��&����������9�L��B6
�8-��A2�����.nG���_e�����.�)�W������ף�
��Y�&��)��Q~O��I���+�!���f�P��+<�N��P[<��DDZ��$y&�{��e�
eZ�"caI
 �4�zf=k�	o*�+�X��㙘�W�؏6c j��S�4dҳ���0�=b,�ԖF-�\M�=�pU�TO���l-&I��1���*�][	���vd�]�@�z߻��*����^p�g�>Tn_8��֗AK��c�+b�&���(�{�l��䝈��b`#�i�w
�����_�W���D�X�����]��۔��������_�89���ɩ�B,
������3�5�/ļ��B�
�u�EouF��������{h� ��!L�7c!��c�Loo �ekm���p��C KF�ȥ�o<�lo����Z`�c�lH��1z�3��3��rj����_��Rr��(���3�?d�9�7��k�&��#��%R۝�1���x
�-�����*�a��z�<�;����v~ޏ�e\���V�
��������$T"&��2zB�V�bs-E�������c�f������s�f��b������]�a9T�mT���r�al.�f[@4!'��E��C:KT��QA���`u�E1wIf���R��{N�ro�;_,��b���㾎^�d9�)�_�<ӯ+)�g:W���F.������A-�f�pJ$��,g��9��#�D*���0A�w���2��[��U�6HנҔ()6�c��F���̾�a�-�1JX-���U}�6����g�Ȩh�T�O� ��%���b,D��r߈�b�XZ�kBvW������e�6��=�[Go��H������B�c`��>G<���uѼ�*�������jY����W)Bv�����0��j��}>�u�Z�SpH��S�O���G�7wd��6\i�#�h5�l��j��z�r�+���:�HS��gvWT��3���P� �����9A�ϳb)+�9��q�+��U�^���>'U�9d����}A� -C������K����/O�-������Ґ3�Qf�ɚi�U�kRSprz�8��]��3����p܃��tU�پ!��b��DpSq5�U�2arqs0C�a���-�̇Q��m%��ա��4UO��H�%�w��k�Md�
v��t���_�N��~���\Ap�M ��qu7Q��L�VA�x֊��PC2��͖g��6qV0�Zo��<ԃ�(��?�(!ec�턋9��iBf�b���u=�nt�� �0�j�͔����!�
�pc��g�H��R�>�S�  x����a�ȣϳ�6�aĹ�z�x)l��=.���Z���k9+����_֟;�7�_�G��d��~��ރ�Ip7�>�k?��|V}�`P�Q�a����]4N1 ����o=
+@i����ܮ�f�ZS�஺��4K] ������N��W�bZ���|��	��~�Y�]@�oY���ϖ��������a���I�R�����o۸�1'��`5m��*7ŏ
9�{B�P6�1a���VA��&Ռ,���u2`����X:�\����3�4�.�gT� �=��E��F���V��󮯅m�P�ݎ<�X�n�҅�Ύ��%+<J2=qǭYo�/�HW�jH*�Huנ(qT�h�u3�g�L-��l�ۏ����tp�|F=���qK�W������g2!H���2��ͭ��<dd>R�Cي]2�v<�d��~��Q�/���0��^���N[����H����l�a�Ks�E��-Ө��uH�OD�>�Z�(p�o��m��0ybj��Ő`���&��ZyFIѢ)�-1�3:�z��H���ڌ>w9瞫V�]4A:*�B�,�ۙ��q��J|� �mҩ�,w�q��I9��Z���h������_/�~n� X��ӏ��dYx(�X�Y�FQ_�"R
�w�u�'EL����"VӢ�+^W�wS���E�5��c��a�8P��r�E�>�"8���GcF
2_ �GVnL>�t]a-�x��=d�Y�rS0��$��L���iT��ă�H10)�N;�g�}�a�=���b�F�؉����&1:��Ä��E�9A	�S����6�T����
����2�T���^��=f����F���#�VՏ�Q`1�N�0�G�|*�9y����ɬ�����r�w5�m�v��o��M��x}���U��>���B����s��&q�B&��03�"%�%q��|����CJ�ަ��v�;�����3�=O��D6�#�$�N$�+0ɨ� d�o����c��K�)7��0z��þ����X��VI�,� ��Y?�Ǵ��mI�Y�.��:�Ax7d���1���ɇ���V��c�NxЇ�CO�%N݁XN�
�"��pX��asr%��u���D�j����ϋX�fڑQ�� �X�#�s�֓C�g�F[i�s'�־f�jǧ�f�����}X.}�x�<o<��C�7�S�'^������۽�c��er�IF|�4��\�ώ)YX2A�i)�db���rr�1��|Nbc�Y����|o�U�0֍��Pl�?���)@~��}fe�4z��B�J˯�%]m�L�_vGP��N��\�����O����� ���%܈W%
�.��v�[���쏂��Fmͩ��9d/���Wz�B� �E��G�ϭ�r\�t.��r�*ًd���)w�m�[��c�'9`r*&�pbt}���R2��zȸ�챊�m �c��l���A�*�ynO1׆U"lB_g'׼ĳ�mP����:��Ԕ�	^���#:�k��~�<Lr� yOhr��h�=�7aG�|^��C|BN춣݁|�QP�c4�N��X�[�GP���{�<E���7��כFu�s#C>J7���j�Z=�¡�M>���\��	;� F���+� P�m���i��r����i�g�s�Y�!��>���n�U�<�~FP��2I�a�ڍX�2+����D.}DWA�}�/
�4|�\"y�	x��/�/���5~zk���t����xx��]���&1 \�쎒��)�~�ju5N�+
��_�'�%Y���C�&iFM���M������>0�,`������L�vD��lNVh���WTw{j�J�G4G�.Ġ��:C��s�Q��z'WL@�����F��+���T�Fp��m�=�K��Γ��r&�7V$��%U��������q7�6"�ڏ�4�#�`@�����5핦���cj�a`����Ԅ'/`���KF<�bVD+���e-`��:禳~G:�9ܔ9�~�3Y��k�g�F������)M��L��0{�V���دo�	���	`�7�{��P���}�l|���%����,�ηjg���xgJ;��:Z�	�+��$��*.~!�J0�t�,�������T��I�ۭoyR���NoEѬ�~Q�1>Hx�e�	��~�WN��lóZ��Ѿ�����p�Ł�p�m/�I�[Ȁ6�8$��9Vi�Z�,E۴�����j�ȸ_� "��P��t�:���>S����#����ۈ ^I��cj������#�l�xO���!l��9�,�â��0���SQG��#�		�V�	R�	�r��	u|��c'���l�f�9�*�1�>��L�+3��r������q;�\{|��Ly{^u&���c��g�kn�����-��KR*�c�_e�!�@�!�7�S���^��S� ��uC�b���{�/�
�R�h�Z��S�Ӭ^�����5�gD#X�Qi�Fp	�i�G����/�����:���{rj�7W	,������n���Y�;(.�����fv8��?���w�:��e��<w��O�d�n������[���/T�+�~]��!{y��(p?.^f�U�g#rŐ� �OVbBP��r����t�cP5�.XV��fkn��D���ʺF���.d,0�jq�;ܔ�L}s����Y �"ʴW���,"y��T�@,zյ��v��Ɗ��)��dZ�+e2�
[����:;���$4uy�M�64t�ٽ��Ey�e��%�,9ݑN��G�.��<qV�����i�|�_)�����V/�D3��S)�,�!�e���-%�y �W�G�':v��!nP�W���7GЁ9؅���S�g"(k�2��@~�F�����!S�j����1��Ґs�C���;-oD��#,�53f�(]��~4!4!l�B����B�z���'Б�QW�-l_oĐ�%ה5z�ȁ֑�A��T(#��=B� ���Wi��,_�0��(���[ae��6Ax=�;����ǿ��A�1f)��k�
BKN7#{����;������+�k ۦu����c�o���w�	��t�1�~MNv�î=���-�g��MB����sE�%o>�D���7(�&�¶�+��Q��>��Y"G��&����XI��	��|�.��6
�d�q�MdH��*	�%��SuBiN@����c��x�Oj�E�`�Gʨ�Ey�6�@�@��q��XY&p#�r�L�Z���h�qGy�q�}fj�᝙�{��n�w�W��[�',��xtK�.�Ok�ˮ�G��a�R�>F�\J��I��ju�e� o�8�F�E����3��7ET��	�A7�ހ�fX|X\Y�<�o��,��ܥ@\����xA�	�S��{vq��5�zj���Hi)�r������@��7�Ň;�M|�g�Ay̶���%t?x��|o\ѥ��ڲg{HC�|]�N�~�+�\��ib�S��8�{sV��l�c��jP����/V�/�-%���C�v�$��x���7�,�5��F��s-Q@��T�O $�--N7�Iú;ݻ˸B��m.ۋX�4�+0����:��E��\���rjVgNr���"����{���]kr��fh��]���y���6��{(�ٚ���T������t�`H�<C�#MQ d��H�}����p�ݗI�L�%��">���p���U" �PB�����b�-c4��aa2��f�* <�y63��Uğz(��(�Q�!:�Ԍ�v�fc܇?ܛ�v�4��2�Q�k��ٍΏ_	�/ֵq���8�ށ�gîy�M��!_�`c�~�/����RZ��b��̤��H�@�~K�:��.�~����[qLާ�x�h��J�L�� >�W��q����=��o[��ػ�YM�拨`��E��j��w,���wP|5k�7(����3�L�o�m�K�����|�E>T,���!�[��T�	�*p�>�4����-��nW[5��k�3�kc?��<�-:�fv�W�̳=����?���Tշ�_�χ�駾!́SR���^��m�}4���
����e�u��Hb+Ω	{����䟺��BQ�2�F�^w 89�a0e8�h�� l�4WJ0V ���I�ت�	���g��#LX,��^ae)A��K;���&�С��/o7J(~La{oO<-�X��P���GV����,������W�����p+����
�mK��n[��^g���fU(�@�o:^:zʺM�X��t�b-+SK=W-��ڒC�I=�ę���� �g��7ڬo�z�ں�=�t �S'j� ��U+1o�p@��ǜlsl\v���e�>����>��=�ǵ�SgO��,H���F��A^[������]�F�;f^���9��I�o��#<��R���d��������^a�""�
@mPn'�w���TQw�n]���D�Y��hً-�N6D �^��ű�J�lu\�i7J�ȷ�i���K���5f@*^],��N|]Z�uAA_����0w�I|���I��%�w���Q�wXl�'��nBiw5��#��KZ�yf�v���p��2�F�A�=<�H��{�<�
D�E���z��an��V6%�lh1>�%�8����0�]ԙ��'Hp	�����V�� �_��w+[>�;{=%;��6�'h"*V&�p!G8ϯ���U%�HS�s��5	R|~���'�8�J��R��f�jW٧���j��10���r��D\)c�em}��e��#?Eo�*D��,	\@#���$i[\c��e7".�ӛ���2^�/����i��)�aA�J *�	����q�LC`\O�_a%�¹�Sf����H�@:�Q<���%�}W�'O�P47�%3>�hY"�|�!?ǨR�4p��t/�
�������;�N���$L��_{0*U��Qu�TB�_6���$XV�d7�0n��`9t{�)����~�Q����&�r|V��J�Z��>J/9\�d�I�I���C�D�������b�o��U����������KYpF��r��0��z���_"��Ő�-�J|Au��x��cb�T��)�����YT�7��hf0H��cR���c��J_�si(�P<���W�b�C� -Y%ǯ5s�\>�A#�C|f]��I�P�l}��۳��LK���j�x�v��%Y�x��������o�\�!,��}m�Y>	v�b��fqn�EO'�d���8����q�;�� ����KV ��u�Ř�����	c��G�/��σ��q��F?��>j�A��b�w*�M���(����3���nfد�>K##ʝ�Z�%3��3��&%UVB�T'W)��
�X�&��y��)�樴�˺ p}Q�c:���*�����֜3J�u�P$
���f�s��'�1mN��.�@�o���6�J�W�cqɘ$�/�T% �t�*�e;p|���~��¯� �#���ٲ^��M~>��l1���7��7�����I@����J���>�fbٝ�]��������o8�/�IH�t]��:;#�K��CGܹjZ�� ,�y���X�����T}2	��Q�)*���U;Ղ��z���l���
��9���d�j|���H�2 "m��aV�;��{�Xj���>!	W�.q�㝔���/#ykRE�T��� R��W�#��e��SB~O'ݳort^%��;{�0~� �����'ZU��-o��`����Yƅ��Q)�>��(�(����w[Kq;y�'�7���e��}�$10\2m�B,�CtKR����k�d�x����,}�
h͞�yMw�d4�p�Ye("j'���e!zЛ!���]x'��^�uv`iW\��5��#�(a��fI�T��k��e��w鰟O��	�I�{p�k\A}��[��k�$�me�^Z&W�cO��x��M����U�}d���e'ID׺�]�ӳ
�|�[+��<��
�ʈ�ϖ#Asop?se��"��]�7�����.9�6�i\���Ŷ��E�h�wj���v��#2Z)T������lT-j&"���Û��q��fY���(�B�����{�������O(��hr��`ܩq�R��N���CU��o[E�����R!5X&^�l{j2�����o�����*-mX���+�G|���ŕ��q���1ڹ�t `
�1H��v�y�rY�*��<�����]�?�^U�~ŏ	��E�_a�Y�w
<���C�h\O��n2,FC[lK������K%X� E.�N�s�g�Ɲ�.��폤�cA��?�+v�~��V�vw�%��QC�ā�
KI��s�oM�����x�6�5��_�c�i�*t/f#��cu�%�״��ƧTb��~[���6����D/P��O���b��2�_���5���9ǆ��퐰]��<`�u���[*/�T}_���eU�T�����%辮���������7�� T��p3�+�)XMEE����������[�+b61e,:E�vb�{�J�����Y�������Q����	�jḿL�DH���o�i�w_�V$��=`(1h��3eJ���N�*1�(��V�a�=��W䳉b��^�X]S�W���m�`s��s�Y�u���B�`�'�$�p�CC�z�?pY��FI�׋d˗orf
NF0�A�M��{��������R���}
�D����ۉ�]�������9����5�0���M��O�tsB5�kF�V��af!�u�������:���/\y�PRF_ۓ�W�vI�۠����qJ��t+����@lL며e	�1�x�#&�52��{�5|ʹ�G8���J�2)��	ZZհ;���W�gҽ�I�6���b�3�Y���>�s�2B��$" �>�N�.����9G��g,�x�ZSP��H*~*&�7F�8=�(U2�Q;��0��|�W��$��Dާaq>O�=��cZt>�B�&t�Y�@�4>:	�i�s	��A/�Î��jF�v:7��v��5�[�#�A�dC̋Y]��=��(u#/�������x8�rGS}������	�O�m$\�Ez�c.$DLε1��!�q��PA�T>E~��^j��	��1��d�*:W+�)�����b�����NN�p��T�[ʕ>�-99ٛ_0��_�Â�(.*�?��P�Cxĩ��n����D��?9\�G��f�
pi�(�<� ��|�P	p
B�dT:X]�^O��T���)+i�<#�/l����e�f�r����1{��iR�h�;�ė#G<����3�U�����#(�i3=�ѭZ���E-z���	�_Z �[�g�ke�����|���3t\�
Y˪�Q�-�FKj�
)���r�G�0hY�����`��"	!d��=����M�2� �}<%����"Fwb��p�O������kxqo�c����Ә�Qc^����F�c��x+����G���|,�v��݈�|�j��t�J�/bK��n\�)����e�Q�����evf� `@�Ɖ�����O�������&�w�9�S�*�68�Z��I�v@P�]���@����ֶ�Q�Fd��&�X�?�ǁ���Թ�ַ�tg �!��(@����/�u�&ҭ��0
�fQ�u�&{��)[��!3���h��AP_8�-��GE|{����ϱh�X��W3=���6^���6SF��^��3�7;��Nf�V�&�'0�[��ַ�<H��8	ﱈ�OV����,yQ�1k,����Z�;���V�79���֚4����wCKGp�jr��|���ΐ#��^�ʉz��?�,�s��ML� ��Q,+r�E�7�"�	��Z ��lNH�A:c��4.�?�ԥ���`��d�A 2� M�����v�_��J�o�b�H�������xmXP��M��-��Ձ�X�� wGNä�\@,ڐ"Z~���3������������nB�^���L6/ tL6+D�n�� K?�<i8�F�x'����.��(��v�}%�w}�}�%�5E@Й9HgM�G�[h�nO$����������3f�ש�J]��"�_� �+`��{��$��_,�QC����'N@=���1��gۦD��T�Mi�W1�1/����	�}�e��N�(��?��
t�Y���h�����i�Y�5��&�)�p��[�"
2򕒑Y�Q%McDaM ��"�sf�[E<*3�r���:R���8=x:��ہ�^�!ª=�:7Y�OV����Hdu�WԽu���dĹ0�ꋱ���Q���)`�[����/�|�:���e�*K�=9C?�~���	�8���5pw���d���i�XBNP���MV$pʗ�堘��8wqy�{`fl�-K���/g!T���(���";���s~��/��#-t�/��/���i+��A!�_����RM�,���&����7�IzA�>7 ��e>fƆ4E^�OZ�i�� ]9X{s��/��@�#�y@]	.B��Ж�NطHG�Nh6��V�E��9�iY�ԁH0w���^�p�wV��p\W���j�!
�j�bh8I���;x%ď� ��3)Ъ[!�4�U���C�.�dl:Q|B5-s�k�;��=� 	��g�ƻ�'G�T���,$��j_@�"*�Ǆ��ٷ�Uio��-�*���ѐ��bT�D'E{k�4
���j�7G�6�A�#���\�'S��{���bn�խg�xr���{>��q���@1��Β����W��q%�o)�Fc&��O6��)�L2<�	'�7�e_���뽛��?V�u:�o�u��|�vxM�t�f+���l��$��d�vI`}c y������8��l�zJ� ��di�;��V9���|�Ǽj����}w_*�vey	���[-u6Q²��pD8ݑ5
'��X��=v)��W�鈽p}{��L�8R$f��&�kw�{o<���婨�9CvvygUq^#��_$��"�f�<9��W�@��<%Ҳ������ϔ�:�ͧ�Yǧ��?���.,�*(YUNm�L>��i!ȡ<��MPN�j�ӄ���d��I8^ZVF�����)w0��2��7](,���o};ss�J������ˋ0r���lg��#'ڹ�4f|Oܖ��K�z�F����fGўydQAP02o��|R�h�����������Pc�9�������3lЗ���X����7'vU�"�~b��/F7�j�|����4֫6�`W���m�׆fNо{%�AĚ�,�����@MAw�v1�Q|��h��CT�T����Mk	s\rKw`s��p�P_ĵ�3�8�\�oQͲd���G<���%K@j�x��q��Y��$�az
��K�W��n�#�[&����T5he�{;spz1�vŪ��L���n�Ć��T��˅�����(Wo�`'�1A��\$�X,�-i ib<P9/���/�(���/̴&��Y�f����>(�O�o���u�F�)@�>DT�:�a?��Q�G�uB����' ���B4��y�OL��rx�����{X�ق�@��j�y��LP�
(���{��f�;D�gG�g��xU��D��_�ȏ>��R37Rzv�@/���}>]���f�[Us����@�85/��s��%�P�$�:v���NCW�T�/P*π���l����=u��g���m���Rj`���'�Bi[4�����]�a���^Z�PV]�g�T3_�w'a�Ȕi��W���Nv&\�� �6ĉL�ƽA,�&%��Ϊ�K��b��8�B4��l[�};:�]e?�S��)z`_Cwl�/���4��l�Z4���zZc�@.j���%�z��ۊt�@-�͏�])��#*����ٞʍD]�"�H�b�|%1�t)�Tn"�[]$���  �*�����p-�d��ӡ��{�-�|�n���� ��7F�p'�k���B�fU~�e���DC�.M����z��O�at��7}�y��u�vPY���^+oev.��lƼ��
[Q���vT2;�H�(�-���]�֥���/P(�n�_j?T���o�6$Z�'��./ ���ʫ%H��>�8�MV-�(�(v��F^�]0)q�s�~z=t ����(y��zrũ�9�w��(��$���2�J�������>���Go�|yP�C��B�<�-σ�Ix��RQɣy�5�S���MlY���o�j��DIϭ8B>>7�x�BP?'�l��
T��54Yn�	�_&�d�ĪOn������N굓%�Pk�{��ltw��[]�U8�����Y�rRE�3�<�}ӱ��Iop��~4��78�a���i��z+$�#���=�ebdT�04�eMU��뙳��(م~"U����_e��O�=N��B�#�8O^kA���0�-Y�#�#��g��m=�����S�6#[Q\p���[ڵ6�ejO^4�[ׂ"����Y�1��0���v��h�i�/H�@N'�l�#�6�MgN㞆�s��O�]�UM�[��	 ����̨���.c��Ƌ��w������NQ��V�So��J�����b��;�4��
�z���6{-5�����J�Z����ױ��lQ�&��	k@��xG��������As�Bi�W}I�ޱC4:��`�-sg}X������jp��lEj�R��V�bu�&SD��FqW8��������U�;PR�cV �ڌ�£#&ɒ�s��I����W;N7�cS<h��|�f=A�ޙ���uï�eF?���{"�)/a�m�:	>t?���&��k����3�bgXc��{N�슅q8gZ/���̇�}�.
����k^�Q�^�P}��H]�� �]@�z����k��K��v��O�&�S�`\_ �nf-J��:���03���$;f�RpL���I:9�*�}��b~���� �`��ˈ��
��nOǝ��F�Xӕɚ#�x+�͙�lhB�������ۚ* p�q�����2��-�ݢ�%����߇�2��=<�9�)`�*Q���a�{T�>��'u0/��+0�縌}G�)�t�X�(�m6�k��뾪�EM.��pc��\vAd�N�A������u�7�7�I��B� �3޲.Цk7T�	��)'|����	���q��r<Z`�AHt��wI�����y�ᘯ(���^�h/���j��"�;z¼+��\P��ѾE �r!�e&t�����%�F
�
��^@'�=���NRB浥*�QX���U�yx�Vۆ�@� �7�}0�l��M1��w��<*q+�H��b��l�����1� *PK�S꧜ڈ��We�ChZ��||P���[��cz�b�2p���D_W���ac|`(�e��_KM*�r��2��������!ȏR�3 �y��Q�%�!\Ɵ'�.G>$f�%/��+#��RË����Dn��@��O2$}!�r��Ŋ�qK��`lr�{�0��������[w6ڃ/���������π�']�Y-�F��֠<�U�d���G��Ez�S����G6la<�I�}YUg��lO���:}2PQb��"�v�)�@T�"�jV�cq7_����;o�쥊��np,'k��s�� ��l#Q��J�rګ�,�Ev�Q6���p�c� ����'kd�p"E����/\<���/9R�����H����'��E�ْ�9�R����(Uբ�'�9<d<�gؓ���R���_��%-��"O�tݣ����\�ƅ�ڲk0�>Q3%k\V��k�T'��X�E���ix�!P�q}E9�:5�_p��Ԁ6���c��ch����Bsw���3W�-�͎ЯII� ��F�b:}�����-|+�]x*A
���(��q���[n��/]�</�OSU�uƱK�;n�y���Y��u�����+V�C�N kM�BeY�8�
��z��j�C@̏��_�*W��ƎY�Nq��B����_�,�JK;¿�Mkן_R-�^5?*[�ے�D*�%��o��oS�*<u_o�M<"~����Lh���v��h���]��\�)b��\�'z9�� � O`g	].�����!-�%�$#ڿ��-\s�q}e���ٓ:�L�Nm����3Oe�D�~n� ���C����6�#e�oBz;	>��O��M�g��Ơ+�F��Jg;-�\d�<���?7�5?��ړ,*iҭ\���7!_�+��ϟ��!ܽ�����i��`��Y��Ya�L�(��J���ރ*�ޭ��IJL��[_"���#�PI!��ί$r b�
i�+�����| �ⓦ���R�P�=�?h�j�p�Y����2(_�,Á��z�:=���͜^-M�����Q����S<���`ʺ�1�� �x�A@E�"`�'��jP�d��5�]ټ�[�>ќ�4��g`�q�U��A�nۛ��g'f)Čj��JyDNY�>\#�0U��TbNK��	��n����ꜿ��qZÌ
5`2<&؊\�1iF̷����L���kg�h��'��Xgu��nHG�g9"�I���L5�b�5�o��̙�O�*EP �~���	K�;ܐ�+ZCN�ؚuhᔑs������R/�A0-ܣ�>���L���0�j��Cf��SpӶ�eA�D�Y�"�����U�
�6��V���+���=P�`ʬݽ%v����ERE-�Y�\�D�5�o��j�\�fh=_�+�5ޢ�+z���ʬ�e5����p}�����E�@�}8�@yå�ū_ʵ��4���P~��S����g��x髨�����	�
���^0���q	[&�]�,7���l����sa��"$�U3q.�k��5V�<�➶Q"��~��1��fG�O�زm��2��lԙ{�W��ت�g�f���1�����Vf�_��待7�_�D}U��V��q:�2w����t�+���� ���a�A0��X��ڎ ����ll�ԏQfH�� �`N�����&>��ؠ�-�|{áE�~�@����tM��!t�w���L����,���zϏgT
`��E�9tF9�x~tRT���RxK��*����o�G@j�Stɺ����l��V����С���,)6��; n��8�� k� /8|��%�I(Ş�q��hY:�q�\�-�����L�v��d+Q�^��[��q�k��0�MWnI��'/D�����Ay�)�4YbV���~�e�Vy�o|�EB]D{Lj�AiG��n���"l�p���&A`)��KyA({/��a��6 ����/�Dˌ���tėU�5V����&�k��!&�e�|����x��	���}�+~2}I��L�kOd�>�lF�E
�z�j��d�x/a2�7%�2�[�-z�����7���BT�h�lK(<8��I�,�PN������%dbA6ƿ+���AW���@~x��⩯��P�&�a�#�C�\�Ig*-)^q�����R)V�:��ktx;B�W�=��ڂ6b�A	|L5!���dGp~֠6[��L�p"A]Z[Y�l��L�[dZVۚ���׆��Y�	6��'�)��'�~��d��M���be�&�-̎}���2��Zpm7��5�ٖ\*�7�ʁ���r�z��,�Ӳ%L��)c��������l�.��oj�LA�z_.��nEm�'�6SG���Z9a���c��xF�
T�W3����)�'+G]~�*��J�\�#o���y$r[*�b�>�TX��ε�pL�bFc�ëo��1�f�����Hk���~@��Ϧ��������xI�]}̤S���죇^C��F6���>�������g�޶�j��y�Ԋ��%����
7���©����V�f�r��;��w�$:����͛�q-�NY#\K�f��BS����r����iY�Ȯ&��eEr�����%=b^NB��(̆��!m(��P[�j�fj�h�$��a0٭��a�\g\�U�n��Jߛ�������A���vrWY�sj+�Ƽ���O�yB{*��|M�%3!��-��6��L�r|v������z��#�$�y��Qts����%_���3m\�oqk�j�S�;L�?�5�l=����W*���,Җ*SƗ=t�w��
�d#@`\f���H�x�+�$�_fƌU��e_!yļ�X���.O���-�`~��DYah!W2���Xj��W�}�uٴ��u9{�8�{����t�V:�Ϧ$�F�~5Ԝtm>I�l�a!fWq�:�(�ch���") G��G���r���i.+nH(�����-�r��Ϣ(&��xX�c�UC�y����T|a?�x (��@��QWt���n�Ʈ������(pJ���)��@zo�$�����K?|�R�e�zn�5S��!|�f���5n�v����q@��쫂A#��q�e��"J6%Dqؐ
�K��"m�s���A����4$,���&X����b7%�6A��i�s��05��z37`��Jvjh�����#���a4��Kd�ߨ��\O�xW�Q}+$%��*{a�?��]�{�OE:#���b��?"Ӳl��~Ҝ$7�^��ʋ��D�+�vawp�����R�a2u��f�U�yQzQ�Ҥ��5G$�.�/��FL7�L�=̟���7�8o�PރT1f��D��lt{�{�7��4Pv����&�,�2*d�(��n��֬F&\'�jw� �ޚW�����˝���c��KL�US܃�
�Z�������YPڜ��}��#1��@vU�!7d�4`bL->q%�pe>�Md���Y�B��-�9�ʦ����fsV����Nw䅍���3��UF�4(�S�X˪�f/�I���Ig��I�e�7��}�i��]#���l�+j��[�I4����8����a�9t㪗Q���If�K���P8`�R�#l)J�8�����0F�	�dn�c�(3#�܍58B�;?�7z�|H��ٺB��+>x��9�,!�ǉ����OH��^+w��G}�,W��d���X�Y|�hB�U�3D̕7{;;�[X�z���ʺ�g��<,�{7gb[���~��Bt��{��A���:!��~��S��6�t��hx�|F	W)��#�g��<!��tbxN�T��!��@�����[M_B��� ����׏�h)�b�j1�@��+�u�A!��'�.��/&�3�����Gn2�����,�G���Fg���n��M9����K�&�������x��W���mG"䤱D{��e�喾��L׾ٿ{|��ͅ�O����*'�=�X���|5ۦ!p�����
�u���|�L�2׃r��ΑO�?K��Sw �������^=)qQ���
���rݷ�J�`�Y������Fuݐ ��	*�3Eϙ�,��<��i�K0���nþP�(�����1L�(���ёi�o&���
�Ҕ��S`ePv�S����ٚ��qK�`�p�U�)�"c��y�D�9�?�Ar�;��������5�'���ԯ4P��(��Be��#����+��i�9�h5ا?�(�,��>���#ע/@����Q9x�њ�N,	���c�ဌC�*k�ٽ�ꚶ£1+��z�0��V~�"
�
F��#ᕝ��_γ䓓��f��-����.��3R��ox��	��-[ͲV٧d���wq��O��QV���V�3�<:3��!���>���י�'[Ǽ�y8i�������K���=PD`���o��t�Rej)Oq��׾8G���hv��^�i��V)��^�#��f�vV�&v���ji�cj��27��ܱ�� .���I1�|᳌D`���1#3���P��f����Pm�E�S�vʪ��C��	�yM�
�S�؞�WU��ͮOό-W�sm���w� Y#g<�ț+�Bs
��y�q+M,�7[궧��1��wx[�l��Gjۊټ��Vu��9��+4�R�z���I�pY��
���z�T������	5����v�c�)��ݫ�����=�:��XꤘY>��T������q$�G�O���<&��	��A�(߰��S(B��~�{�u���QU)�0 o.:���8��/v2#�l�{���\�
9x Hԭ��Z�Lv�>�A�}�0���6�}K�@���l����y�b���v��(���A�L���-J��7�<�Vo�k��o��l�dD �����<�������|� ���ͽ�M�gqͦ�� ��n�� ��-�@`�t�-�}�4|�G�b�o�:��~Ϟ�?���ܷW�6���h-ݤ���X�J����f|/kZ#6�*���[�e>M��_cyI1I3�3��<j�����06�}6��Y�N����Dđ�|6e�5�#ѝY��4Ł뵵,����.�)_���!�4V�Sƞb(��͊��Ӊ�������_`&wCk�i!Z�䡹%O:<-�+�n��xI����0�}��[�_��}[���DJ7�4��>#�����9�ӎL�,^L5j^�-u<i�E�c�u�n'������2Ԧ� tIuc}�Ns^
x����D~|��궼�@&r��m�M˴�p�b�^�7��q������%�5��0�7i�7��(�	���A����$��gn���V����җ9���@��5���dp垴	�ߖ���z*I㉽%e���#
W\��8j���~[MT�A/W�tڠ����̒V�ح7f���9���j=Pϕna��	+�b�Q�+_;[F�^~G�%*�4���,�S5r� �N�q�_��B�+����^KR���4>��~�����Γ-��;�r�[���g5�3����D��!��[Ҽ���.J�u`�^��U� ���J�D:����"�LΙ��	1���c5j�!�6�h�<��)u y<�9K̇�Ds��o��I��2v@9���~w����'���Y)�����N�OĬ!�J�9��Z�C�O�H��Z^�+��k�Ҥܪ#�����BK��$V�����Eg�I����fݱ�F���Q��-��KpN��O�i�#�����]���H��O!�&`y&�˒���ݫ�D҉�V�gF<�,X�n�2�7V)g���.b]��K�⏡�$]Z�j
E�1p��� `we�	�[k���a�I�3\.E���2R�����[2JS�N���4_�Ff|&��O�*S���S[V�J�T�>*�hsp.,�Ê�K���ԛj��K3a� R~ #��G�J�Ry��|��n*Dz�;23q��O`�.��U���p�X:>s��Q�p7/��M���i��:��>{eU�@��*�Xݚ�}��]�A�\�&����(qZ5^�����V�F��i0s�s2e�}��ǦZ�ߛ|���A��8���G���
S��E�Z#��~
q~��*Wْ�7�;��drA�a��j���g���|�����e�衊�9Q��켉��v}�4��ɯ.�=�Ade ���C�N�݇�t/<��ɲ�0��DB��+��A�^\�}/�����p��"1[��i�R���:`1P�~K�m��:Z�0��o��X&�����o&N.��t@�]V�\����02�Sԥx�(��p�i��1j����Ak4uz��f�O�t8Λ��jt�����z �<֕��~a�3qM�O���C��ßrB<�8��V�Խ}��r��7����G�A?���K�e3C_?����m�d�`(kHVX=�!:���<���v�:ݠ&�={ �ы�%��v�/�P�tV�;%ғ5��c��c��\�y�rV���~e�c��1����CW�_����QMw��{Q�p_���Ͳ8Lل����~����Y*�h���d�$H3�$��,&�ѥ�NS�_N��Ôږ�g@���S�>Z�ًN��L���$��m�l!���yM�<n*��3��Fv�׮{=�㡫���w�^#[�e:�0��K��\��TzO0�Ի�'��s#�jt�z���b|�T���B|s͞.O�L*�i >���J&��oz��-�C�r��l���*M��~���_�+o�&oU�n�J��^�|���m
K�7�R�c�BM�`��<vU+A�Yu�+�J������]�9�8���.��1z�'�K�F����� �q~��W�]<5���ǹ�ĥM�е��P�c�F�*<J�b����^�������P���5�L�dQ��#�QP�X�E��_<Gi�R<���H��7�G�I�6��ĒQB��㫝� ьr%X4e"�d#�J�UM���"AW��`�:1�3�ƃB`F{x1�|t���*���]�Yv9Voy-Oo�Cũtm���y��TKI7�UV�t�\��	�oBY��j�{ �1�%z�%@؜���|�g+���0�Q��xu�w�x�Z�r,^�o�ӯ��$@�}`q�r62�5�e�fl�����+�r�19�>�>*fa��,�jMCg�J;�_Z@�'ܪ�T}0R�=0�pZ��z�&u��+>R���a�\���	����˳$y�h�P��H �M�F���d+O������� ��w5�qTI�O�6�� Jr�8��8��3\��gX|�=�� ��RT�`w��xGZ�� >w~��h-��4����&~e� �5%�����u8��Q<�'��OQѪ~��~���|��c�?͌�;1A���w;�!1�.L!m����C��s,b�QJ�ʝ�Pq��ZB��q����|z��Cg�ȃ~1jB,Uz��7j	���U=��/�N���8��E��3��N�*�*m��M�'�k9k�Gvթ%|ے&}Lg�<�	:�V;�L��Isd�C� ��cL�;��v	85@9�#��������~g+֑H�
Z�0�1&��G��A��Q�t�d��,K��"�c��Y4$�tz�Y���Dɱ�+�[<�4Et���w���k��["���(/h0�IGW����#G�*R ��lNwt�u�@���?B�쯀D#9��0�q���r�o\Ͼ��(�cc�?8�����P���I`�5m�d�t"b�}�hZ��)�t���3+R�Zx��;��53Z=c�"asA��L&�������S��Y.I|ɫJ�Sa)��j�����=�<�lF䟧�7�N�:��)O��Շ��s]�2U�pGn������9�wJ��}������\�蝖�hsq������e.w��UѢ�D����1E牔᭿q��X�+��m��ajf7ʱ���`���=��۟:����g�SNs7S����1W��hʢ���qQ�J��]�,А�f��+��AwN~~,_}W�㐩�é�&���~�����51u㰞��軣�)"ˋ��B�3����. +�o�I�iމN��x���C|r˹:�S��}Vݧ�~m��F���P��6I`/eV�.��] �w!"8uO�!���pc�<�\Q�5_D.�%�D�e]j�W�@�-&7ߝ���CZ=�����6'Y"�x>�JN��]`�,�}���WI��~��K%<=��b�[&Ӊ�y�G�o6]*���.b�"��j��ϙcksg�y�klk�DWPR%*�`����c]��V��|�ء;����͢\#�a0��Kp���s���?�e���|�{�ZƫǍ_?�����}$k���t�4������'��<���A���%b��+KB�c��'�9��1�P�Ƞ�~([?GOarF<��a�N��N�z�k���$��JW��(���UH�=�������W��	p��$�q�~ǜh�9�"�5tP�e�CޛD��{�'];�r�*��+�Qߤ�Od���q�Rv�5�vf
���h8��N�ec,�[x�� =��ץ�2������\�ls�G�k�fˮb��o�4�F��CE#۳gX�iD�ɺ���(Lv�� ~xM�䱹ޠ�-5;��2��v]9��ן�SNq�c��'U]�IH L/
(^h��d�\$��m�;;���~+�<�8́����oG5 ��}ߤרQ[suQ IO����L��[p�����D���%��dxȉap;;���F�g��N"�Χ�'OA��C(�=uwv���$��E��Jza���^��{��1��>fFg���N*�{P�H�*
�� �H��vَ�FYR�lYVy�"�X��{Vh�Ձ�ֈ��Q(<��n�1jp!�w?	�Y7>?kET�h�p*]����&"Ptے�_~!zΚz@�<��.	����'��|Wv���E�(�o}G�~��&���=�ι9�zw�qG;���B�$~c	���	&"`�)�*����w��򳭞0 m��"��Dj�ý[B`�+}�F]S`uw!�L�{�8"�%Ԩ��꩐|�Է�+9@��j�6f���k�XB:F ���IvO��G&�oQVN�H���M�]�Z�4��տӦo%�\ +k� �	H�&>4��r6uh�)�I���؉�?��!�$(vRM[��[@8��-.�'�A�����j=g����l0�����������2�I'��)ac?�ϴ*�_���\->T{p�&�����_�5d�6�v��	#�$�r��M���H���^��;M4Ge$3��	��Pz+7��E01�a�H	>�Y�Z9	���:�"��*���ۆ�q��ټ�	W���{k�H-�)�7��X��Z����i�ٰkR��5x2_lp��g���B?6�ң�CI[��^,�.����݁ L�,�Z�wbu���q�ų����.��c����b�k�D��M�m�-�1S6���I5��<xڅ�9˔�*��r���v6օ#]�t�#�%��qG��ȭm�`s�(�(Kyn³��+��_]��C��FR�F�v`�m����HC�_3�z)x�u��Dk��}x��*^�ӷp9h��I{e֍6�Z;F�O�
63�jڳ�i�h��t��r_i�u���g\^V�l� ��C3Bޟg�H&f I����N�&x�9�E��T��#�<b��H���`���6�v�-VU���Bo�:��ϩ�x��hMp�T7����F��ctE�E�h���Ko|�X��?��%��f�>��|������b��^Ln\�I�<����m\�D�_ץ�(����#2	u|
�i�$\H��"q�� ����[3{��.t_2��@\��l³L� +
w �K�z��<���pw�J$ᖲu����
*�
&�-�Y�����=�<�mA=��D�o��(����N�1=�X��Ur�=�����N�c����`. #Y��
9'Y3՘��~1��i���t"���-�7Z~�r�q�~~��<����]�с�4��Nق3g2�-�|���I���)�6&簛�U�+����F;�빸#�Q^`$&$[a_̡^�$�5��{x�g��j�`r1G�"+S`0��m,�{)E$?K,?�Ꭾ�4V�yiK2daŁ�%�]���@�xg��U�(l�̕pVQ9h��R�K���`Ƶ�跟]x��Z��
�������h�'�b`�@_�EG�j=�X7Ç"��;�Zǘ֢�D7t��I��������YJ��f�r�&�b��K`�RN��I�m�n��l~^�y��e;�u�PꇃH�z]�c(����n���'�Pչ_���o�R'��2�q�\��߃�>#)cH�!���NmO+W�(�'��.�P_Sf�q��2��
vw^�&��/����<i����c{Sk��,����:�Q���3������1t�tY���KQ���p�)�����XىBԠ39��Ht�v����I}�q-����BP����Bo�^"nƆ.�o1�E�uzk��]�"WMگ<�G��i�ͱpř�8}�73t_7�ڛpyjИ����B1�dS�B�H�X�\�,kʈP��uб�����c�k,L��2f?GE�^����T6q�/�+�ɨ�.v�"��@x���'Kr<�sۥ����?����髁)����`q�Q�Ѭ
E�U�лV��B����V�ԅ�����e@�1�cG����Tbi��5��6*�������h<}6J��0G)�x��?���RR��p2��f��KY)�9-H��(�OIH(�eB΁i�lڕ�����l{��I�3_�HhJ�(�"^o�xF���T��H�T�����-wQ�ht`�ˤk��{U}w��H�64A'L�ļd-߿o�נ�i��t�0��LA�tfK:��ا �8��Q/"�~.�x������;K�XЦ��m�q��33R!��LV�˰2z�x��ʤ6ͳ�Kl[�B�AK�L�����J����o�| �:/+��LQV�c�5�<`�uy�!��$7Ea�k���r��S"���J��*5�_����!� !�OU�����6�Z0��1T�^�,�\#i��m!�)� ����D:���]�6����tN��𘓛�=�(>��:�0嶹��!�Q�x%�J�,Oj�d=Mn�Iuj��)��qv�0������(�{��S{�������c+J�;�m��-H��_�.��:c�W�'B�f*���0{_�B��Z��M�;:ޚ8s���$�&�D�������m�5��0�#G^�2=�6 =بr�x� �#��~����xO��Ҩ����_�ƞ��:�y��,$�@J�DFQt?��Zt��_ॅ�<���ة���\6%���ȿ(���=�ɴ��^֣ �jAN��[��� #�)���л�^�Ry���1I|����C3��(�&��ﴲ���{������ȃC5��d�23y�=���YZl�BmV�@@L���G� j�E���M�S�o�E�r�dN�n���|�,��YK�s����`Qe��F"�E� f%���:X��ah�]#�>`A��p�v~���y��Oev�A�X���8�s����º��8�N�����ozK+Â���z���2ud�,���?L�JY�=�L���A�P8a�&�QQ4�0|l��#"�y�D�:@��Q\f���=�j��v�8󠆲;
Ȁ����3q�1�ت���єr �Y�����XY�6��M�x2��[��e�ڔW��ȇ\Ɯ(�P��,��֒=�?,�����?7�ڮU�`%�;�T�U�_ԘLmc�Z7���#p2z�vE����������,m��SziNT"��9�S|�l ��?��S;���[ȧ��W9s+Faڻ���^ڴ�e�ǿX��>�I��=mmЎ"����ϕ6�0�`�0�E߂@�X���0����{1��}YnƟL�r�~}�ۉ��yϝ�H �j_[`�H���4J]�cNf-�:�*XV���w�s�?� ��m���,��r��r�:�,���:���l���_A�J�J��	��)&��G�ަ�Bvp�NڅU-:1V��������āxUe�R�wI[z�G��4Y� _uc�׫5�9��o�sw#l�� n�s��~RB駀O�k� ��7��k̎c&��=sѻ�2&2������F�/�ޙ�����b�~\Ip�,�oz�L��><G|X�`[�G�A.��`u���^$s�L1�>yD�,��j'.�Cp,{�[�p��G1�s��>v�o�gx����Pe�鷇s�:��m����Z�4��;5h~�JuH��b!�����Ż*�:�$�@���Ζd<��k	��p/~���ʴ<'W�']^����P�4l�I0�#�dh�GaL7���-���N�����v˯lA͟0B�.�.�j����W�H'e]~�R��\���{��؀A��m���Ю��'�Qrm�Q���<�Yv��.
���2�;�7�{�=�e#)��	\��)seF	:x=��:`B0�T�v/�G�*&j˨��Y(��'���� �)�@��/�s��S���I������謀fP��ݏ^n���,>w(4ZN�p���ח;��MK7A�s�c50S�ёv�H��߽ވ Y�<U�: ����Պ���G�ߡ���"��6u�rF���*})'Ɓ�#أE��gNA\B�C�q0|:9Ik'��+��gt�id}���?d��<�+��܎��;��Ԅ`�kk����[�y�hD��P��N3�	�[DNJ��}P�����Jd�v�������-a��9(5��;�ԏ>�DnԨ�:�+E�V�S�[�7��������
Ej����V2��̵(H��0�y;y��l�L�|����������EDo��O���Ŗ��cm�e@�_"��=��́[�����t#@�y<�$�߂͹��ښ�\���E�"U��P'��J��(�ga����u@�7���s�EM�n?�A)���F��~T�|�T����O���	�*��@�ι֗^؅_>�XV���|��,�廌��P}�h�Enj,���e��~Hug |���f�Pw\�sʊO��V�с9�~vR0�곏B=�tO�HC��!����w�����[��2EI��F>����uG��NA�|�9d�Jq+�����/5\�sq��Ay����v�>"�����Hcޔ��W�E����6��CTԶ�<�[��D�lz]��b�g�z�~��b���	!�w\hm|T���uMl�uf������2� 5�F;:��C�+��{[]9�~4ԏ0�xo�|��X��܀(�g�̅�_KЀ���	 ���E��/ݱB`�twa��Ɂ̈�FB�TnA�b���`�	�޹4B-TE�� ��;Kԥh?z�-z��f�R�@h�F��T�Fl>�'�܂���Gǜo�^�{�SǊ�ȴN���S]�q_M�π�u7]J^��y<�jS�J �}u��o�WK�rRf�2`}�f�<E.yۅTX���]���p ~g�ؤc�c�<�į��D�-���}Qd��譇Z����QB���lHn�H��WFԔ�;}�c�$��Qۻ�`��Y�J�*��8k-�X��ܫ��&Ui�_�TZ�&�i���GmY��Ѿ�u9[ؓR�a}��B�hLxO�0j� l�N�d�W�H*>u��a\C�q�P)O��
�8u�չ犛h/�)�t�r@����4�oi��ß�~]�������mV~���?#����,��k/́c����F:�9�����V3Q�~sʹ6���F��y!�Z<L��Ǐ�̏Ո!-h�e�ǲ"z2���6��_0:��d�!�x �i�^���B|v-��	�Ȼ}��w\��q�;��䊇�t��Z�g=�^|��<��`����<��gWq["9��0������-yw�Ex�cD�ԉ9��"��?�_��~��i�9��奮]
Z:kp�e��zz��R+��'��������݈Wn�H��(�Y���8�eZg[��~Z�&�u@��d/Y���הPn4� ��F��p�V�.NB.��0�idB�b�;ݨ|e.if�����Ƥ�?Fo���O�7?��������߱��U��D7,1�� �̦�Ԗ�����j��ɂ3�D��h�FZ�. ���Ά��m|�V����tn��p��E<��P�"6�5��p�J�X#��Tζ{���B�[j��Q�3�A�gU]�1H�C�h0a�煖;99 �/4��:�$$���wo��g���٘�2҅@��������� G��
.F��?�%`��F���e:-?+p�*��Tg����#�}U�$�u-n5�,�M�Ie�Ҙ�ݺl?]R��*�̿P�4-� ��;T>��ڷ����
�������o����JF`z0��.����oY�}��/������cV���)�\�u�3�����������@�B�q���x���0Sc���Hqr�CJ��Zq�<!1FS�"iXm�I����M4(��������Z2ߞx�M���e@���������q����u$C
mY�c.@cFL��	<�V������t�H���@-��Ux@ �zt�z���pn��:B=�U�M푷*w�,zU�S��bXIC�V��J�a%�m2@�+ͺ��!~��]=q������in(yyg'�EC��h@#�$�Ixo��uF��V��o�s2��������F0�@d�v�Ek�iD�zՌ���X5��2�g�r��[
�> p2��:��+�����9�MNW�����Z��TZA.#ް{��5$ ��e�{���cе��=��w�mU�o
�BɛD�[t�����. =o�|��Ʒ�r�kt��f`����@KP�x��{ռ�Շ�9�#��9H���c��F��5����b>�-1ݾ.\h?����Ŋ�m#R���3��q΀f{n��@<����b��=;��zU�~ xd���,�+�u��cĽC�n�0�5��Ⱥul\�m���?u�l�gw�"(*ª�&�s
k��M%�T�qg�~��=���ɷ�b4F��/s���K���d���N ��!7���v' ���İ���E�Ú�[0?U����:�CՇ2&3�n��9f�"�Z}_�c҈����F�o_Y	���G�ڤ����d0�NԴ�"���9$�%?�n	_��.ىU�¶��sB�>�%�T!vp
�R�hD1�V�޿&Jύ��鹚����l��C���O�%��J�^fL�&����z�_j��"�'��~,/L���#��Y�Isʖѝɥ��j=��=���l�Fb[ߏ���m��-@
��uoa03k�!���2<+
ɼ�\���.u�~`mLwC?!-��H,ݜ�+��w��+���$���i�((��@�"�s�.���+��'�3}9D]}��S��-N��/=�ÔT�oK?�Z1���0�!�A��ѹ�h`B0Fω��(��{�����Y�@0�v�s���Cty ��n�ί�04OGY�Ca����5��8���zEKSI���Bj��m�q�� �O�ʕ~?f�U��8�͚�D��������2Z��WHG�O�J��!��)j�Pv��?��F��R箵h�����%�5,� C�]rA���\��� [ i�� s��qt��f��ml�+v5��X�2�3@��te�������.>m����$�巏nџ�Eb��(#��l���j�f�H[��/�6��<ğ��xoQ�pn���h1:Y��Ň>��F�n�j��D�����ָǷ�NL�V���:Q�'f�����[��pرI���9�o�cm�~��W(y�l8_5��c�B8�.C�g}z��0x^����(dJ���\��N�H0�¥�4V 咒�m�;��I��͚G��
�}j~�����u,�)���Fo�'�0�:d�H3q!	0���9�ӿ�%�|�@�V��ݙ�a)�j�Z�O� �]K�"p��n���/����w�4<Gx\�P�ߨ��g�}��s�K颜�P�yqK-)L�y? �� ��]RAh������rV��L~�Ʃ(��z�8-�ܦ����	�B0r4��8�������j+�0d�2�>o�[ͫy#C��;#�Ҷz68��#y)�@�U�Eб>�4k�E1ey��/�y���0��R5
�4d/�N�7�����-�1W�9���N�j�X�\�?��a�eIǻ�B�i8��3�W�C�e�ݢ�n��|�(�hWP6s�_41�b��Ȣ"�\��-m^�&����������DM�������7@]E�#=��͡,���z�˾��B�V�ބ��!�	-�;c�М����1� bK��:�c��8H�7���G#�[F8\�|c�������b�� ]�Ncf�1ƍ�NE�.?�-D������y��0����Bʊ~�j����X� �N�H_6��f��;�[���.�,����5��Yݥf����#��b����L���	DzP�ֽ����Ү��,e��Y(Ҝ	��[��Ӷ�e%�tW��J���r���2Q�W��|�>�GI��Ը�A��{�x=I�)�KE�/iN0���t`����4.�a�U0��1)��O�)�B<ܲ /��i]�y�>�
҃<�[.�Ӌ�G�6]r?ȩ"Dp�N���3�L/�q�G}�Nd]�*�Ή��J�zJl^���N�SO݉l���b�2�2(��J��o�/(��I2
#��c���%N����Sp�ȧ3Xg�jfo��R��Mt���"F�dS�?����@@����{��Џ�n�Y�E߿i!��N�*��:"�-��� ���H�O^���kA�	�\Ճx�nvX�:~���^n��<���
z�?W*����i~˸0>4_"�'�X�=�* y#��
6�e�,��#�g��2U��Z-�U�>���U�����������Ro��+މBS2}�K��5�C���?lc]�Fm��Ed2#��v�vјZ��|�ļ"���BYY��-d����G�%�=������IS��Gs�%��"C.��:c}d��]�ɚ�2X�S���}]�&A*��en{p�Jq��z̸e�;�5��ԙT�L;���:� �r�E��V >_;���p)<u�aF�1�V�'��uj'x�,��O�ŉ;���Q��F6n�����Ğ h�: Ɓ�Ł���0z�S
>7�CU .�v�����I�Z���{}��Y1f�_�ܔ�~%�U�q!�,'�v���w��o����Ze
fs�jk[���~L�)+>�|�FtArU�<f��{����2U+2�z~�R�p"�_�@'��K��qh ���hg�/Q6ab �\�Đt������W��*lO��^�ƷJ�#�39 �"�X~�N���纷���9���d��'{f�������x��Q�;>���ƛ9�����G䟵T6��9H���V��4.���6㮦9��6ADT�ݦ P	z���=��)�p�<�d�#�a�{�sP�K�z�j6s�1JkM�d2X�^@�S��!��hٜy�,�N���+�yw�tθe?���Dnyļ��R1�e�^�H�!��^O�����BEm������L�h-Uז�S[R����~&�+2��;)~kŲ�F�T#��m���e���<�N@K�*�6�F�Ա��/ןÄN.�묠?���$������w<��}jCщ5*�$�h�
�#�e՛�������O%|�7�4�`1��R���c���A&u��h���*]SSt!���1��_�������1%Su%�HPXkH���va�&R�������~��h/��ڪ�.kt�OA���L֖t��B
yd��"�h����*�:�%F�=�f���a�o�T�I��v�  ��q������������v!9�jd]ƩE��ǳ��:] �6.N2�yG����6Y���,��7Cf�}��{= ״*b��1��7�A4=yW��:ރ¦B,ZU����r��u����m�3����2��<�p@h�
���L��x~�]#m��6�q���3{���S.����h��_k�T�˥ࠫV��������S�(��0���Y�u�Z҈�8,�YD ,�%Ϋ�`��۲�Y�����#�)���B�@f=�?a岺̇�<2G�Q��`�b�<�)�-$�ό[~<�l��Ԝ=x.)a
��L��6��j���kBɌsh�k��z��7y�;g"9��qR�G�:�aw�	�XT tT��'�Ӌ��i�[$8+G���<[��Lh}5 Ci�tL���D�s�NU����-[��L�,kL?��I�[.Rsܚ]�g3H����,�Qթ뿄���D	�vr�jf� �V,��Dh����^��@�OhE /Y���E��r��*z�I�ͦ���?�G�n��EJT�gGρ��f�0�{�"�O�l�`Zsʞ��O3N�_?�HiR�ϊ����K�5���*XYU��lu�4<�,�C'\�����˚�3��&}�;��r!�sJ��STi����f�����&�9u;j笫���� >bي]z$�ve�l��X�r+w����T����b���+A����]G�J�J]�������*dHmJ��S�2��ze%,�y��^j��*Q4�������"�H��t��d������w
Ҷ�r���	�#�&(,M��c�=�ڈ���w�_��<0��(
��QM�%m����Nɗ~/4�FqᱢBd�9z�T3�����)^8u����[o<Ś�nK=&G����\f��;.�zd|h�� [��9�Y����X_9�;�����m��H��*A��;�l�Y�|�Wq�Z%�0��j_?�Xu2~�3�ۼ���mU�&E��'�5�lesL� ���-�sy�.Bԉ��Ƽ1�N��Zv\��sK%�,?�f�`��cb�R��gQ#Ɨ�0G�}:o�5a��d$��(�[��y�3�5�J3����}������wj8c�ņ?ތ����'!OE'�B��3��ٹ�y�A��%0�^ʹ�O�[�y�Z���>	,������#O�� ��D�n0aH������L�ֆ!5�-��Sl���w	X��'���?�Q���ܶ�p����4c�*.�=+�$N�]�4���PN�����_*vZ������7�C㌷��p@~�F�̍	e����6����z�̇�ځԂ�&����h��Y r���Z٧^����:�L~���>���
jA�J�f�����TX]o.�8�&��$(�&��B���	'�W���r#R+m7�;S��w8Z�79|���ߧ��#S���?/F�N)w!��Za�r\��I� �y��]x=�.>ޫ�Rc!I�nD/U�G�ȸZ��������j
E�"��lg�s%_���1�K<34=��D~UY�%�	����K��Ƕ96��i�U始b�o�NH���Q���GЩ�.|���*�ؓ�Qw/t�	6�;����M�g����n8!���Ж�`��ʤ"�	�C�@9���ۤ:��s��B/Ff��M�<e��4	�߰~To��@4]a�R8�r��x�.� DU�ivT�?�W:m��'}���Mx�YK�3���n���ɂfL�. S8-f׊��H{��*�,��kr�z�'��2H,r�uG	E���̜;&\cH�&�����{*�_�#qA����
n���Eh[eW�{�ֹ�Lgk�"�՚*42B
3��d�'�3���m~�֩:�i1PD%�2���Z%t%r�7v<�/o��T <l�J���A��5��:`�>oD�s0���Mü϶�|؟�����$P��(�{�!֜���g���}�%-B�c�N�I����H��cB@C(X��()Ur���
���R�t��<-L,����!����geec�Q|U�J]UsLH��N厐��ظ��oh�?:iQ���'�λP�P�8��^O)3E~O�5fio��8+��Q�jez���V��-��W�0�¸E昆�[0{�_׏r.d�� ��$Ƣ*ǧ������qEuE/�2�2xӫF�n6��y#�})����(�tI�	����R�vT:�w7'�<���q0K^����0-W� ��nx�˔�����W��fO_@�!c���ʍ����!l:����;}{trX�>�(3��{�	��$�&�d���-�0���-U	*��j�EǷ�68a��MQ7�e;�w�N]�^�^��+48.�UJ��..��D�R�yt0�޺�`���d�OKs����M;��b�3;�ڠ�f�k(�-ؒ<�|�����fA~��*�;�}�i����0���Wp��#Y�8qwCC"5��r���郞���|�[W�0nT3� ��P��^�a���+%���|o1h/���A3zE�h3,S��n wQf��L��F[A�I{�t�;�<!I-���8�jʬ<WE��0p��+]�E�E	s�bC_60-�r�Dd7�!� P���b��:G�#\F��k�D�\D'���ԫ���zuo�ޯ�ф�꽂����r�U�{�RZFR �"�w{ՙ2������V���X�1�h��z?o9�y�kE����z���@`dS_-DԂrߔ>���{�dt�]w�x����ȯr�v*��AN;��@�#�b��'i<	�a��M��3��r�=�1kE�8�5�N�FwS5�%T��9���\h�˩tm�ist���G��k�_G�Wo�j���:l�W�u2	K�PY�%�Lr=6'ݡ*��Z�*tՒ��Q���=?Q�4�ӥ�
ӆ�K��;�o%���ؚ�A����t���lq�V��U�`��$�����c��c0#g��ɰ!��̀�!���EH��i�<[�t{~��� �?�����5o!�I%2F�u��/�`�5������0e�K��#��xC;����}e����T������i$4��Տ�۫3"=x-\}��5���LC���H]z�4�	�FAs�\Q��>	�YwR��V��{?�GM�@F��{�>�\`��:+9ϰ��C)�Tt�d�&��2���u�p�ru�����5\Fȡ��.9�r��'�����NWR�i/U�>A<^L#�J�K*��O�3&~Aɏ��͈/Y�`g�Y�~��ؠ��sՐ����M��O�iX��:��Vfu��H:�����X�����c3�H����� �y_�52��Ccrja'��y[�D90�Šac����(��M�~x_�����:˕�k�������0CO�I~���ءU���H������;�օ��R�j;V<�x�V����|j���eՄ�#���}�	�(+���V�A�Ԍ��M�5̙/@M
��F+��C��
�GM'�`U�0C����W'�䱸7A�ГJ����dڄ����x�`l̴�R]����sX�-�Rm1!��whv�dD��e��
� �%�s���H:!�!�X#V�y�&�pQ�ھ2s��XjUU|���޸�-'Ap���o�q��w�
���Tb�	&c2� "i���"ϭ�LE�N�-����س*�;�8��4P�n�`jJ� X���=��td���?6;ƃe[��8��b�D�m����Pʵ�'��'k�e���	s� .h�%5�'�1��Ш��U.��MA1��c3)��X.�_�c�	�q��}�D�T�Ki ֑�2A<7�}�OjfbO��Ca�9쬓'�׏�7n�����!��`�%ط��'p=W)Y^���9RL%�y�J�\թ��y %���k�[�*���:j%5��+5�����gQ���7�T�X!O�_��`�W,=wX<���	�R
��pϔr�^��R��Ț�Iuold�ұ��|G�g����f�j)�m��~N��e:+l��rvt�J��t���Eu�

����pv�4|?���~���Q�妳��#;-�U�)�kg}NU�D�>L�QD}LC(\��ٜ��._�FC�?68�A��V\j��1�G��In�~,���El)���3<��I�`M�����x���ܞ�R�<��G"�ʾ�< r�ev�>_����'�ǵ	�i?�Z�Օ��4��\��(�[r��S��ï���*	Q�s���8�*����Y�e_��2���@H�(���RMe8NU'���&E D,/g
,�p����ư<�?��P=�aO�o�f:4_����g��L��i8p�`F �t"�����	3�����yb��h�f��h,�!�e��SC磮8(�cO��ӨN�c&�!��������I�	�uk�B��_
��8�%%X
�r�:���P��[T����R��
�qg��[D|v7����+)����H�a���]����qX�*\�[��UO�4�5~K��v`�m���zL�zAH�|�G�j�i� h�w����&�%���+R/���Bjt�k
x_
k�%�5����e$f�F�g�Ky���8ĵV6�l}�u$N���<:�Z����&�s���m����εk�oG@=]�u�ar�]���*�Փ�KПM]��RJ�m=3���X�6~�WԠv#��tM�H�v�h'*|�eT�k\�ֹ������i�?��ܹ�(-���A�/~�4V��~�r��h���ƚЯ�l�Uy$�� +�<@�4��^!T�k��^�Q�xƀ��%�)��T����Z��WC�r�ZP��	~(�Ԭʅ�ۚ9��7U�^�+-*S���u۩�r�w}zDG�$W���i�k��%uX#	����of�A}�~�[��L;'�p�G�^��4��;�e���̊��$Ӻ4}q�GI�=��C� A�l n2�n���0�;_1V�������4TaqJ�T!�xJ���s[]*��R�F��c�[��a���O*��n��5�_1���!�iA:=��Fb"sXCR��u,@{��	I��Fw��������QG�5nզ�*�xk��H�d�r	#1���+�N5�&�٤�}�`p�n�d�0��%Q�n��{���`��Q=T��Lr�۶��C7��=/�҃�뜻e�ΎՖk�;��L�NɃ�޾�t�v����	�����BR~2K@��&)V�?��V"Mp�s\q����aI�?�l ''Kã��N�ü�0G���|��u�7=W��Q5�KN� h����Q��[�w&W]]�E����b��ɜ��?���}���B�W&�wO����X��^�VH�ʢ ���-����=]��V�ȩ�Xq����3iY�!��6ڂ�cUzaA^X�]����8���C��>����QM֚�ȼk��a�R�k=��=�<�>����8�S FU$��-E<ۜ���K8� �z���5J����B���n^6�݆���?��s3?�����	���2�pZ.�Z:�N�S����O��V��@s�]C�Y���N:�9�=3)�g�&4��]_��]9 �Ugw⛇��+
HV���p݋��7~z�����g:㰒�{b�0f������.b/�+�_��ݶq��)Ҩ%Ah����+���<�j��L�������R���K�2����xgm�����)��/��dsI�'�$�"�sS�-֦�����k�xV��E�!�./C�)�6B�d��M�z���	X�" MMb>%_ϗ�H^b��?��~|������ᖧle�l��'>V�&v����d�t����i+��>�S:?�h��=����$Zm���?>���k��m�D���@~�fW���lJn''���X� ��_�]����%��»��R夒���0�����[ߒ+�U�":�m]��^��Ix��6ozdgl��()���,���v�n��0�-��}�儌�ԃόb0 5�]!wRy+F��}P��KHV�;�m�&�#G���-���t�[v���$�	0�4d"՘z��^�<KSi��{R]�ISeR����zؓu�V��kׂy����#��6�+���Xɞ�����21�,����+�o���̳Ƚq��}�L�6Lwբ����$IҲV�v��.b Z�"���j��X�]{]��%x�i>���<�tB��q�
�e^nFL??�%��2��Zu��W�Kv��]�1Մ%U�wT�k��)�,0�n����l�T�	u�k�Ģ�U*D�5G_��}=�d���� uUR�5S-��)�c����I���4W��U�c��qAg�Y�4X�b&��|�	^v`0Y&�uAh"R9���o��pg��:G�@	��얭�&�0�{b'�޸�#0WܬEٝ�q�d'D}+ov|�=���'0�����#�@.�h|8-�G�7X_�`�X0, ];y���"�(jn�>n��^�}��I�:6}�#��6��&[Y��\���_F��B�P��Ph7�>�eS��g@��	�l�R�+�u�
4��sҥ>��.~)"����܅R�7NʅT�L������t���'�}�6t�%SWF���v��k�Q�����5�e��E5[^�.P?7���r̯�����+�`m�pYh�C2u�7�?�WGU�z_֐���?�d��_NNL\��[���EL���ꛬ��B�l-���WhA�_ϻXL� fyE�"u؈�����
[T��v��.~T6u�A\W��C9����'�n>D���e��_f�{�;L�����
2�V��YnL��+n�[�
�w9DYx�� �,Kx`���Լ^^�r|g+�+�ۗBi���2��N�I��%l���ñ���aL�����73����]r�qSI��x�9j1ӻ�' #>��k{p6sF{�K��s8"��W�
��c?�v���������� r)�7�/p��H��rT��ɮ!P��+�4l��Џ�AHu9�j�(��c�ElB-�U\j<EY�>��3��f3�|��Wn���(cH��Ch�t�)��`�#a IbԤ���5�R!�^��4���-uk.ǲt���!����*����],`�ԐT�y�w���FU��z�b%��^��7�y��Wc#��␘�z��I��a��l|��pvI���`w���A�N(�3������{ ��y�}{�Y$��T�H�����1��<8ry�Jz}\�)G���z+�v�f��0�<�c�Sdxw��&�tp��,;V;�'���U�fSՊNz.���\|�<�ݤ ��:��vo�+ƨɻ.1��\�}�Ỷ�!���0��Jg���Ge���[��#_�t�(tc�0эfkٝ����N@c��ܱ���}3��ԟ���
���i�l��; iE�:�f�Q�2j���k�/�N�a]��c���h�VI�@�P�Tar}�z7�X�9��źP���'�r"a�O�E���S����B�wc�I�����l���}n	��"�S�׼g_��8h٭}��x�ĺWID�}�H�<�&�c h��ʉ6�^ǱV�v��_i��q^'_E¦�Sm�7����=Ӣ��o%cl@dX��&�Է#ƛ�%F!iGP�}�Ym̒%������Ε�%�7܁k�5 n;vr,��E����7�@����f���*���y�Z��`\�`�Ѝl��И��dgb��,�R��JT�  �=@��U�Y���u��2S��;���+w���e�3� >cD%~��Q}�P�ۜ�6zJ{����^��];�3��0=o?K�s��N��$�y�ȪҺC����{S�z������~��z�[u%K�T��!Fn��Yr�*+�<�n���h!N{�V��Ҍ�0��Hfp{��2�u�Q]�\b���'�S$,�C��`�d���}Rt835ǁB�I%]��Pa=���( be^�w�A�Li�`Wϊ:^#4����M���@2ï,�)E�9	$��,̒8
�� 6ӊ�4���bpT@������W�ĩ�Y��R��0#���I��@�π G8U��(������֎�⍬�dR�����{8�o�a�,��s��c�kh"y�0���8�s;(;�򙸦;�#L�X��,0y%a��F�hl\�I�^��'b�j*S�Y$u4�e&J�����Ա��A��<r>�DO�?�uP"X���;a��[cF�Av~T^#�b������Ȏ�ثB��(#v[�X�Ze+�E�B?PR�V�Zw��@_�5��C&å�,iy�vR�NC'?l�P�h�*�SI�P/�C`ˁ�dƐq쾯�H��|'��Zc;6��KF]�V|Q�O����|�dH��U�����W��cBx��`�ot% q��.�,N�
(�T�PxJO<)J]䴛���Qά��:����v�\ �%nَw��y���$���r�m���",�ʳ0���E,07�D�L:)����	�GB4������� ��72��}��΃(����*�L�uG?�A�oD�8K�i8�k�(��S�٥�>���Us%��h�08���-�[��ʾ�4�� �f�68?��4�^xW̧.�"�yˤ�e�^f�=Z�0[%�� U��D��2i�K����$��L�w�$.z����ӂ�h"i���g0��@�F�������k�\ࠨܹs��.��ߐ�]�-=ȃ�I�����>��>��'
G�;'���(�d�5��y�:�/�;�w����]�>{�bV8Nkthy8I�^^W�=f��V�,�6{�M�~`� ���S�
�j��l�N�Ý���Ia��fM�oSP*x� ���#��]���i����	cu)��P����xc�<�߫g�J����&>Ɠp�cz�<������J��*����.6}� ��N`=�n����%�����ߖ���	Lx�}W��zWp�P�P~�@�q��1����,�ߣ�} ���C��'�!�)��6g��O�|5p�;�ڢ���Ũ�%
�Kg&��*k\���c��:� �_���l��\U2�s�%{s�~n��Y]�.�jۋ�����T�q#o�a�P���I�{��~i�p;)�tD��� :D�����f���ϷO���)V����Y�=�K2IJAԋ��g�Z����_ը`H�@,��%���Y�����=�I��/�Pdh�������˱"��Z�S�c���&��V�zxV��gܘ���bT��>:�o� � ���Fkd����#������R�ǆt[��|�A���]������Y HW��3&����C�r{3���ɞ�L��L��b6�M�C�']b�~v���U\wE��~*�%����42uK\9�֞��p��̄���;��\���?n�.�(i�rJ]�:%�*���9B<-�?�t��u!��y/�d��F7<K<r0i�	��,Ձ�s�*���\�Nh�Q��T�6q[:��[�l\k0�0�����ؑ���!�!Խ
����
h�n9��֙"��c쓛*O���L��-)�^NS|>6s�ų0����k�0=��ڑFO�NOгAj���t�BvI	eM����C:�BL�93uU#dcz�P���n{��q��\����irdf-��)��%�c��ف�	����_��wp�4�pE��p 
1�A�i�N.�N������7��%�ZR�٥-[8�ƞ���;i�FҗL���;\�W^Z�E��
�R�V��LPJy	�w�2�_�?��<�����'5�ƀ�4#DN�T�x���謣5�.������5�ޝ�M���a�y=�)�b��v,�f����G��&�7wy�_�D�c2n����5q���wC�M���_U"/���[�87q>����L7W����D�(5Ƭ>��X4~J$r��@t7��OC>�8:*�b�~3\�S����ytю
���s+�R"��/��{��=��ɮJ_��ޓ����4��;p�Ř�Q�/-���N�Z%�D��'��^��x��`�v���

$���&��.y�vX�M�l���a�[&6�LtZ�r<�����2�Yݬ`5'Sc<�q�����%�`b�&�u EH���x>��l�/��3��^;'c)�>t:�ܙ���,꛺	��h�m�kR�N��>2o�k�)�7C~��=~c��
�o�ű?P�j�����@�"
��hp%���W6�8G
'�G���\�)�dUQ_�Qr�D�m��F���*����f���7z-/�w��}gJh@B0#4K;��3�ɇ�
�/J\���J����TW�҇2��r�rݍ�q:
��Bb�[�,�&
�y���Y��U��6|ei� ,{�g���{^{�f]')�$�mSj��t�h0�ѱe|1����yG_�?o�z;uMMx?��~�y����8Oj��f:+�p��t���㾨d��>�.�K;�g"�N<K�G��U�g�7-B����/Ȟ�eܠD���wh%�B��h$)�鯒]�q�·o�7�<��_���L��-��hH���u�%���2^+�=+�f��[:�2�ܾ����G$l����pG��b�R�.���,���>}����.>�����;G�,n�?>���v;������4��������_ ����UE�*I�(_�K<���屛rc;4rf'�x�y~������_ f"���o�s|u*��~�ڤ�1�wd4ߢ�R�,��:��,�������|�f:�>&���#d*غ�naFO�įS �s���F�r��s�)�*c=L�W
T��"����T2���ׯD��o���49��a�:
,����Tvr��?�D[�;��-`�j��	�p���s�w�"��6��Tf�+?:�J���z�>��"�[n>�X����"����|�s�Q���$�,roH̆s��!1W��^�B��m��l�fUn�]'ɸ��^�z�LoKf�TM{�Ŗ�'}��D��"��;#~��*�1Ty��b˟�P��Ű J���s\mj�r���Ɽ�i�-�EӅA������~�5�ъ2����g* ���K
�n=�㫑��n��΄ͽ��L�:�63{O���ϨqVA�|L~�	������A���������h��94��:�Ql�f��mvyw�x��P^T�"�ְ�G��_
Q�y�63z��.{[�i���'�v<t)9���X�0��`���
��_}�3���!Ɋ��3��e0'��vK,EC� �/��aW�L}�2w��ae��[�=Pz���쒦����oQ��	G���}-�v�������W���NCX7�T �E��2yjǂrO�;#�z�i�2��F����.~�ѹa2�p/��E�<:��ꙹ� >7�_3!+"-G�sCўT�;��e?٬��v���?$K}�m8e��9ua�_W�j7���e�ժ=��E|)�d�b��e�S�
2����YD��.I����X���LQX|b�����-��P$}�SQ�|/}9	�t� ]C�D��	sN�6Mݗ�O!���+U�s�P��F�Ơ�ڐ������z����f�����E��#�W�\&є�� �$1}˂%F�Z^dk�{�3�4�4=����E3���U1|��c��+$���V�笍2hሀ�*g�`��D�����ł�C�F�3����g_}����x5�Ńkp ~���k�wyB�c4�V?�'�n��+�8�5:TT3��d�{PH�ߤa��&��
aG7�RL�Z��j/�ܙ�J��֚n�~寸m��9GB-XX��O9�5g9��͂��n)���u��a��X3�:�͂pL2~DY�0���{.�Z+@ޓ?>��+�Ix���F!�ɡ[ޯ���6������U��>�7�����h{�����y����/�Ә/��-���?1'VXA��r���YV�"Y	����b��M���5�~�B�t���L2ϭJac�Cڵ�|l����$$���������u�_���uk�BY4����b�hed3��Դ�ʙF�B0�%_@��\�����ܧ�i��s��U֤ \6��N6���~��o��iw{��Ci�޴��M_3"��C̕�z���T ^���)K��tz̿G�庄ע�vΥ�U�3}g��Y1'��ZU��$!�5no���W�>���Z���ҾǶ`�絥�5o�h"'2=�Zf4]X�����s��k<L|�>��#�p�����}p������LՖ�W�(��=�.#�[�(1���<2�	��)d�B��2���&�|�+���Sޖ�I��%E���U��l u�x���e[����I��(S!��u�u$�����Ȼ�6F_���/�~A�����[?Z�(�=~#��w����r�A�J�V;�.��߿�,]u���J���t��=�I���5�@�ꏑoc�b9�Sg���FL�P����(63f�q����`5���Ո�Y^�q��{�p�`�s���4�⡗���<;JXV$ z~dkZ���<�H)mapk��МF�[/ˠ9���[�����L�c���U�n�������n~�av�s�Īz�Ƴ���[��]}Y�H�!�m[Y��4�Q cM���z�����D'FŽ'i���@~��|�TQZ�x�ߌ�߃0��������������T0���Iￇ!к����-d((�V������N�~1�>�f��#���Z)�57?
Id��-�fCQء�ﵴo����Ze��b��#X!>�h���$����-+�j�B۰nJy��&wݜC��\3L
�K�z�SV���zS�F�1�~�)P����/�����&h�k6�Ԕ���('=�b�q&q��]��88��ѭ=��f���j�r�k5�����婶�V%��c����7:_3� ��Ig-�M��T�Q�sNC| Da��ͻ�S��K���(�]5�`u�*�N7y2f�Jc9h*�ؔb h��ڔ1қXg]sM�燘  �}4-7c��ŘYZ��aG��?`�D@�޺�˝�y��� �*��TS]=�$�%�����AMB��M��P?�5������e-mN\�</I����`mO&�F�
�b���'��k�MH�[�7ܓ�	��Q^H5;���g�B!���Sz�Z) y��G�A�Խ�2�N^��F¾�L����E��O�Q����.a'�3�5��NrI��h���E�N9��4y	(����|��G����|�4��.P�ѡUЧ�u9��'ߎd�ŏo�U ��no��/�4�	4�$�cE�G�"��O�5� �Qų��fB����%w���5�)�	b'L|�1]���Ɛ��h{��h��j�%Ok�}5$<p=�M����	D�ǯ���/g=�c����	]�5U�V[|��~u��T��gsrP�J2oxV������� �)��8���M��]���Q�U �6ڹ?#H6�Q0�_ˮ�W3�?ӏ�e�1�XU-U����p�a�*�Z�W�)�aO����1se~H4���h��ك�&-�4��#sH�i"�����ͳQy`R?�7����0���p6J��~;m,���\���Wn��Z/[�СҚ̔�e�?{D6�Wb�}������k&kl�5���y�4�?3Y�-&n�-�[c���y�4��ρh+?+��e����s�{DS��b�xS�%]��H�FZ�2MX�{F�����s��i�Ae�d�<:�$�_p�EWZ�b����W��j��N��>�9��=���8�@� Ě2�PQ�96�.������O	��S�H�u�1�l)R)���5;�-��OW �>�D݀��H ��P6��|#Ll�>�Y�%�ƘgQ����������+�a4wQqo0F�P7'f�V?����/^��+�������W��s"�	I?�hTȷ=����}�U�w�c�ӣ6��P���B8s�V�z�c�`�|�ni�Lo3 �X-q<�"1'�^r�@��b7��2~�H�7۩��ܑ�s����!�p�I�$��A��Ǹ����\���d�F����w�7wdFuj��c�3f�1%��_�t�����5�';���1
�+��������ӊE�`�L@���bX����.����? �u�ԃ`de�`�����}���}�|!2����s�G���>��u�J�!�L%CH�Z��=W
!J��H/�ʟ�~���~ctU��s`b�b�=t���Q�?#l��W�B?h��nŒ�;R`chRY��km��U�4�_6�d�jDw�l`�-�LN���%n���Ҧ\���L����RU�t"���!�z��_�rI@�m�&
��A.��r:O�{;�w��D�ɩ,��c���/C:\9�"��SGH$�n_[u%ak���a��Ȕŵ�Eʤ���1�;r�s)U6�pMtp�U5;@��lm�{�<U4��ṷ�(��y!s�}{.��d�m�Ny#�W|ctdbq]I!����)���B(kvT,�l������T�j?C&K �0T~��=�XY�g��C��-2^����ڮ%+�6�{�_�-��
x��+Ǔ�����G�M)V�������V�i^��z<���fF�N�2�B@d��iO�&�h����V�6�P7�b����$�W���q�^Wp�^b��;�'�N��w�a�H�3��z����9�Q�W�97��i�t�+�������K1j"��)�e���H�'3�G��c��8-�jO��x��H�L�;�:]���V�<��>��0u��z,���S-��B�������!�� �E�u�$h�[:��8!Y�=_���E�%Qa�z'弎0K%���ri�l-!�=�%��ʯ��Xܼ���?��-`�]
,��<ML{�k�KsF:m�Z���`r>��=�����.��Qp��������:�hOx���j0X�=�4�jT˩�
�<sǧ���:�l	S0��	���."�Y��6Ҿi�P
NJ�X�䚖�[�0��!3V��[ϫ.IN��Sp�+j�9y	�8�<E���k���M(y�q��`���;GN�R������֠��#������ͯK.1�?�����zJ&��,Nh�&�=�i��C+^ӵ��bR:����]8�=��p�b_�NF�������!_� �Q�ulvu�J/��R������n��̄r!�o�-���䷶0��Qf��V[�T��!;�]�� Z�����A��:s0��	J���/J�1!�_��IإmV2��,G�ͽ52���NS�aځ �H�{����<�	�!�Kfծ��6��3���I(�^����~��{�yR!u�u�V��~�� Zx�����������.t�����՜x�0��X��b�q_��y�H��E��,������V�̖k,�D��#���Ȭ�k
��`�bSit��-*���$a�#;ͰF�'k�F*O@�K�_�������w�1u�%�c��	��;�o���Q�%�)~̵��Ot2�ch2���m�T��x��k������f�g�8���)����߀;��)�E���]2#݄�4�TsS`�o��ܑ�?Q`$�|��}������H��}�ô@c���F���K_�;2���������R;�����677������S"/��r�o�c��	��fh�����h`:^o���\28�Y�jK)�p��%_��]�3u�i�by�#o<L^�K�a�f��J})�L	�+h
���C(^���"�DT�%:��W���6�ȍt���j�`Z��y������h.q:�-2Z�O�mɐX
Ȧm��W��{P]K��Pb~O�k�_�VF��z8؉<g߉?�u����
���F*��sW�v@dy,n�<"��Y4d�0"�����t�g�G�g��8�=|q�&�?���u��a/�`Z&�a`ih�9����BW����sv��A��Z��nbV��
�[ѭ:+e��t���'��8���{��zV7���']ǘ|*)�6?])2��ߣT(�O�^4��j����k�I� ��"qCJ�gm5(�˗9LO2Ǡ����
 ;YxxD��i�`Hf O���,���U�S"v�& 4���ݛ�9m
*���
S�d1�n�3�
�a�q��Ej�ge������.ؙ�||�4(zW��AM"��g�(�q�QY���?�
,@԰��hɧ�%���i۸�vb�J:D&�d2,RBh&+�O��Ϋ��ZһzGa�[�NpaXl�刟��U$$�Ub�M�U��1�9x�W�]���MY���V�|B��K(��c{�^�{8l��ڡM�{���7d��u1����>pH��k�5f=�q|Zj��il�5K��:�OR���:�3����9�,�Lϰ�TRZ�C�(yhNh��`>��GC���[��n��I���YXV�;A�nFRu���#�@V�gXm}�d
j	n�y��E��-@#�o*�u�T̼̫;[�~�֛����GKL�yu�)�M?�	�Ӓ̿���E�>:̾(Jb�#�|:���L�Brb��M4��!B��@�[�O����������k�s雰*u�f`Aw�^2�/���C[B��V�]��(�Mr�����=��@�Up�\M0B\PA-xo�3�vz�Eu2?��&h�?|��|�[�O0-pT$������=�k����q��@v��.��z��gZ�S.��<��Y+�V����X�����>��P ����P�$�4앜��5r��>�Y�S���|���jn�:�l�>��S����noln�:�я O=l�������9֟�����<�sg�g�`q_
� j#�:ķ�����D����2�C��
 ��U.���-�}g�m���A��`�Z\oF�G�<�0$s����փ�F�� n��
�7�Z%�������i����`ØFh  �	L�|�{Lf'T(_�f��Ew�"��O]j���>�̵�����M� ĤZ	�;v���Tb�Q���o\��������znL�j/�9h��בs�+�A�O�T��7儨:��2v�w�{����~�{�|�8"��:�xk�w�x��OD���S>����Uv��V�W{�3[D˰�lO��.��B*ן��6��j�����e�Ifk.�҇Y-ׁ*�"|��u>�'����7�����Z���Gry,�䷴�wxe)��M@B�Gc�;NFTA�&�'���Pܐ^��SF�}�[%RW�gv4ux�EG6�r�N?��h!.�rx࿷5�+0{�Q���+q�.^
�8%��w]��O���~��K4�ƌ�~�D�kj,C�I��H�b�- �M5D��3Z1�NW���C}�qp>^ .�:���%���k ��g�ݓ�oH#�͡OcJ�CI�| ��i��yaE�K��@�K�5T��kxf�?5˦�2�;ذpd���#G�夑`��#V��'W�Z~d��`v|b=E��/���7�$���2����B�su�,���������蘷�=��E��͆@��S�ꍖ(if�T���<�:͗?�=�&khk����e�;x��\�E��;w�o�0��]�u�_Hn����vA�U~o�J$���ߩ�ܜ۹x�KJX��k�&��߯�]k���$	�	��I��.4܊�k}�������Y<�[��{���^3d:�M��*�������>.�[󯵀��K�<�[���CK�����e�3Y��3��kM6�q��-ǈ�|�����aKR��^A+��K9I&F7
p�����rHJ�9�5�����["���o�'U@Б5��.������T&�U�Lt~��G^���e qG#�����r��#����Q���b����By]�j5�p&x�@M(�Ey���0ˡ��$�g�σ:��^xw���	ٯ��Ggb���Ӏ)�&i�����΍��^�����,d>>B�T$��yl¿z<�����C�L���~��?�$�xW/s���	?�p�3moTr�V��h�<g�h`��B��΋틛�L�n{�R�!� �4����sS�V\��"�	%nh_&�a=f�eԀ���N�eƫ-��I��~��DUD�:)�`}�D��趐񤠶��7�F��d�Q��{/:VE_}D�\:�
�M�� J�mIz����s�Ѯ��B_ͭk����(ϭ��s;� !���؏��cԯ�����,KS.�6{zɓ����pB�i�
��2%sh��Ɠ�ǆ���-P���w1:�_�i���'�xT�f|A�2{��]rpj���-�J:u�$���?V���I�ߎ;��Z��\OCE����&�nG�DЦ��>���N-Ѩw�����"�P|����I��&��