��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��l�����f�J�éy7�=7?�w�e���˦��X��(|�EN��:D�*��{-� {���hEې�_�p�P�Fॹ(����ұq���[�A�

��я��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����y�GS�N>L���z2�Իͻo�j���0��@��>V-p&Wbyw��g���6�v���ǘ�	�|�x�O�i9�	KKV+�NQ��fVx�o�l�G���^F���W��
3g��Lw=�ʤ��;���1|�W�"�+�K% �%�c�l9�t�
N���ד�ۖ�p������N\^ �����������\�gG1����^�,�����@��&����f1�ӽ?�E���|����Z��y�]FGgn�Jq�����b%>}n����4t嵺6'e�W�?s"����S WF����_�Pq�/�a�����o�	P��$l)���B#�6�b���,x�,�����8m��?�ME�Y�=�H�6X�)@��,�`+���4����[L��g����O���ŦZB�r��ߧ��S�iQ8Y���-L�;�u��7��U���q�?�ⷯy��c�����r�n��F�'�q��Y��0
��OB/b<�\p�´���F�����p��O�r!��X��mV���6��'4I�?�GljO.����ZfRO"�c2�&����s]2	ŃĀ
V9t� Ii���f��mʪ��^�S�l��9��QCX1��_4�`K¹����'��tq��XQQ.b��kL���8"vgb�m�4���]A�R��;AG��A��mi�*$(���8R`G3�!cid�;)w�}b�D�c�4�Ԓۗ�/�KRe��8ݷ�(!1s��ڰӇQD�ǟ���Dp�}�o��M'I?�˰:�Ԍ?���׼}g2mW�+)l�
n�����6k'٦�V8���#3�n"�h�6�~���:��G95�%����vM������Ӳ�=���Hjzb�D�gUҬm^Sb����-�{�J�5��`�I��Q��$�w�x��Yw^�%��s
|W�SEh��/�!S��!�D����9K��L׀1��L�o܃
�ۜ甓�jH�"r(�l�[oU���%���e__�޶����Ul��ܖ�������/��na	�պ�\2Hb�~�{V���f	��w�u������@�U���Z;1�����F^�#�30]�D��(l׍��t5/��B)���!uOG��$�+L��i_k�FBm�~L���V�\?�\�W�&��q�͗�/]s=$Bn:?+I%s��/��9�]���h��#y���u���5|j���"�����!I�ah�<=o�^:�|˲�<%nf�f���]���ٲ�P�e�� ���2��y�J��T�������=M��G*������ӟ�\�2�H��n6Tm�:�ߺOҊ~�@���@�<��A(����I��ޖ�B���n4��Z�j�Bj~�&D<щ�)/�b�hW�" ��]R��_�����!(cWF"����y����T�R�ZÈ?�Xa��j�i<�2o�����?�6���p�7�f�pY���.�k�Z+N(����)��(������]5�Ome-��!+'��sL�b�����OA�ǅzM��9w���s=�E�߾���p���Y�ΰ߽Ԃٯ7�E�/^9
�2�0���|$$�:�䴾��Xj�@Ӯ��<�MZ �ND)��	2�az]R�ׅ�$=Szl��FUrf{�|_D���h�k�g�"	�ן�aY[�k?+C�Lj���e��G��@���g���|�0�T(.n��v����%��m��~�����)�������9�IѬO������H��v,���h�S��9��O�������/3q(ϻsV�#�qZz�x�������yw�@�o1C��Kok}tV�k�M#Z���K���J>2��n<8����I�M����|A�5�(��Kg<Ħs�����t�!b�\�o�rG�vW"����BA\v0���C��E��N��\z��^���4� ]���3�cb<�F��|ԕ�:!/�j�lZ�N�}n���x�d�3lM��ɆS�����s���O_�[�$,�@!{Qx���E��6����u��
qW�&�A��2��6j*$�t�7�s�ܾ��!�x/��Fc	P�EnB�!���{H�+���������2��Rs	�\*l�l�.�'�4���Ā���O�s�/a>PP������#�����>��"��1�؋	ൺ�m��^/��Q8��T�:S4+�-�'
��>��c�]�@���S��h�}�ef��㲽��<Co��@��U;�T}��E�̕�Nio��}�F���@�5��[}�v�:Om��^W%�v`m����& ~]�C�1�z�� �}jA�����I	HK�� �A�d����@&T�V�rn����,^A�a	u+�w(�sU�����|8��AN��R7R	�J���E}jpܛ�ڭ�,.����\uI@���]cGԆhTB�v_#3�M�@�W���z�s3��;y3&�\P;e] (ܤ���ĳ6/r��o�^A�;V�/�}�ז�`/�by<3�M�팿�t&�B�2�v��.1H���h3j���;�R�K��^�`B`��������9t\���&�nw-���/�_��8q����7�s��ʱ���Zb��H67��ӳ͙�	�-(u@��։��E�i)P�������?��5��������WH���O[��k�F�ɬ�b���iB����(_����ߨuLP����;ٍ]���G`9a?q�����>�D\pgx��!$c�$�]�W��b���'���t�����@	���=��v��	}�Y��X
�`N�P!JwR^ޱ�~��B02@{BV#I9��B�/�`;�`<�9-�tB�u��b�>��y�-PN�@ B�w�ܚ�y���+u�l:׷0�+���vw��L��@T���(N�����t�&W<� �W��E��` ��!qD��h�=?��8�jN���RM�`8b36��ר�tɽ����)oh�w�-��4W6��T`Y(���`)��8��_�[y�y�_T�,*�*hu@/�eY��G/��
�^�0�r���Q��J{�'*\�F���\����|8�/�����oE�y"�>�t�sQ�A�(1�{%�᰷���g�*ɔ,���~�xp"&��[�ř����*��6��N(����ϩ�e��Ι�7�o�*�'`<bA�������/�K�����ɥ:H�3�Jr]�-�ԝ�R�@�`�����\د%�c��e��:�aF��o"�BF�o�=$[�cOڜE n�=��GC/��J<&���5��;�hv�I��[�V݉���W%9�p�&l����g��кͻiTy9wz�n�ј��T��rSU!�vx(UsE�x;��<�ؗ�S<zG�=��l# ��O�jY#��{t3+��4�1��4�;��g(n0I��
�����3`ttӮz+��\��W�7`l'�9o[�[xwH ��|�s	v/����9��¢�(j.�H���xY\�[Y�ע��@�quK���-RP� �[L3̜�>�@������ź�w?�V��"�3�����f.9�l�ExW�� ����g=�zi��-��Љ����tF�H,���_�J�D(�H��넷|Z�?,��d�|�P��|�q���lXIn��K��
��_�/��n����;�RB�G^xb,Д�Y=�[�6�y�:��N �K
�#r,�`l�ᩩfuS&0Fr��/�>MLP���|�uB�z��*�hY�[e�W<�,K	�{�
�X�n����0��\�T�U���7T���0��+�������H�uQG��p�'W�SFP�'�ms؅�0e	~��ԯM|zcTɓ>�,�ع�o�ה���J/��X�N�q�EuʶT*�2'>����/; P���+���7�&���7���E�����.-���I�z��E�{@o��fR���d�4�	{/lD^}_�Z"۲�_�Z%�����f��KҸ8�Yo����αc��Ə�^Jgr܇�صLڰ�O�m@�f�ӳ7 Tb,���vc�Q�T�Wz!zD�Au"���q�S�jfK��1?4�#�o�G1l��6!��4��sv�da�K�?�����[>�izP\��U��"l���Mm��=�F��;�ӂm �ǋB_��A� �@���D������H�rR�%w���4CS�1oxlN��1_B"����V��摜y���O�
N5�<����DQ�E�2�]�{?LE����Ԙ��R!塂Tr.�5y���r�A+��1��ɗ�r��4������d0Y)f��-�[l�ai{�)[���x��NRWI$�:	G���L��}��3�j�=��+V4�@���cO.�|�JE$�aT�ڤU/�6�i׎ߙթ���A�$/��\�7�C`	^s�\)p����rr���I��-_����+Q)�ץ#sb5����Y��{}���ӑ��GYm���~!�1��e�] ��B�������݀�ta-�MP`�s^	?�ȇ_���g�ڴ�w��=�V2!��Y�=��3�*	r�аR}��Wbs����7$�?�*o!b���?2'���)D�qC�>�Ƙ�Z�j��_y�-�Z��\�B)�]���dmg�<�ӻ���!%��%弄��Y�{[�G8�0�=	H�z�1zB�a�f��\5<"��ÂLPu���r�L�,n��CŇZ� ]�v�g��Y(�� p�r������qC)��j1ne��^�O�a�����_%Wo�>��B ˗K����?�B6[�K�iD9�v��O8��}�������V�_cZ���Te�/�����˟��-�=�ŀ"+m�f��2>�|Å���$���$ߗ�a;�D��T+
�~,������k�"��zFu(�T�kj׻r�@ˤj
%�w���nPZ{s�p̛@��Z��v���=n^¹�抍�Yſ�,�إ�}o�$��5�"�d��y���՗�(d�ZXvZ�փ�8ո)6$/|�_�d$������d�۸�W�mGFE����e�(t+y�嚳r���\!s��JUm���乁pEL��d]��5��a�G��O�1\�ln�j[4L�W:$$<�>��"�)Zw�ܪ#U&lIX�X��Hu��}ñ, ��\��^�{݈Qr�?	�j�V�KF��r�I����Z>��N+<�xZ�;ЎM�$�q��s��e��(v'�g#�\c�v6�N;S�x׾ D��%\�T���:9�͚��`#��%�]�v�W��X;g(s`���7B�<\\��~^p��j_u�?����=п���S�M{��`����?�!	��t8@�r@�*��~	{5�1ը�����FB<`Gnc�F�wo��/�M�����s�7��QGC�"�K8�<��&꥛ҲUb����:]aV��	º�n�w��t��:b,�� bccQ�/R��Χ��b-)v��������?MkzX �P%:a�J	#�svI�8 ���7C�$t(��~���@فJ�a���;1�/wBJ��6(f#"��vc�Hs�@��o'��uᖁ��#h�uƤ�@���4��nGo4����$���������2��� ��N�O�����9U�a��_�uP�ț[���\�S���`��d����������;�K���#l��7qu(�Ky%l��W�!OF��K�x�&���s���
��'��>lbI:�ھ�I�&g�{qF�ڐ�)���"e�}$x}�kB�t��(�bf᷿�:7'�m�y)���G��2ҝ����Ѹ�n��� ;DU���#]���L��V�T�E�������-s_=�d{����d�x��o��WQm�R3�l!r�90���@���S���?9���3�F?�?�m���0�>��)��	3("BJ�Ѯk� dv">m��A�.	+����?^-/;�������Q�d����E�F>#;��i�9Փ*,�fZ�/��2`�&��f����6k3G��O6��Y/��N;VhV˩�l��0^Z��5G�ya$JF�e�IΞRW_pR/�W���(�a�C�g]i g�
�j��4��-�U,h��^�OV��C[���?	%^�U}�ɸ_\۽EHI�S�aE:^g'�W]0����y+�m����4>���4]Rph�Zʜ�V*B���vZ}���N܎@&���k�J���4��۪��8���d�:���,��v�\��,�M~(&�u�����߶�N���:ɸX�Rnا������c�Q4�YQ���.�C��Ҏ��ɥ[���q>�jt�R�u����S��N�[.K�[�k
̙��dc�>U^nL���=�?s�ف3x ��c1�vc������8�ъ��ɥ���=�6�FN�|{ڿr�c�&|Tϙ7����\�_yOS��W��
L�$�yT���rga]��;���	V�^ܶ�ap]���wL_�@���q.��j��z�9�n	a�R���&����\CTϟC���I��<�D�Ȑr�_����J����6O��V[g���L
�L�z�Y�d��M�4�s\���� ���ʩ$����pA�͇�˿O�0����	_=�՜�V�on��D�A�S�r/�pl�*��k�Y����-��ޙ#�Y.�������u����yPl�#�_C�%�%��~Yп�$�1�A�G�4��{|x���cr�u�l����b�ҳ��F�0���户�o|to��5�T_�tΕ�Ԅ�B�#:fq�ʙ���0��]��Vի&��8n�Z��t�f�^���L�eR��1�S�'����uI�ЪM���7q�'D\K��ڻ>�e�w?�Юc�{c�3vT6.�}ޔ�w�ڍ�NAb�o��:��ۜeg0�=#�$�N\�,�l*/h���|��<bs*�H3��p�veFP��y8T ����#����K��jy�K���[�|���2{�Ǥ�VV���rA���Dn���}hcH��U�U�t��KL �R�aS�/'\�XC��LF�t�boqNs�^�8l��T\�|�`��GH��/�+R����cD3W��+�%��]��
�˫��	� �ǎi����*�U\~�.4�����]�8ig��K���x���U4|���ƕ#��8���*b=U���'�F%G��ѧ�Ɵ�yE��2�Z<���	�F��Ë��I7q�E��$�04�~,�{�պ�r��_�z؇2k󯹾Ϗ~AhhR!�ٗAŞB�C������>ಈ/�k���k�׻��P4�oSL��j~I��S1�{?��<)|�)��؏k�����yb8�4b����@�a`�'\��!��s$�Y񧳱H#�WS�Y3_Ӓt���2�.��A�8Ժ ��ێf�����K��;#���P'C֍�ݤb�͠�g��������SIf~q������h��6�"�� /����}!���&О.����>�Ԥ�=�޽p�2䎘�B4�f\=��]��J�\k`�cC�*��9���x�f����!��,�j�*����P�$��6�M�{ō�v��i�BwI�񘼷��(���F����߮}Y�N&>,O(Y��.!��o�u�qV�>y�UU�?8Z�h�h�SF�P@޵
�_�A����"��ecVl:+��BtbH	7�dH؅a����N�Ud�HzM�*r���~�;~r�W��m�����I�.p9�Qb#,�g�=b�\��c_��V�����I���GZ*o���D��:��eH� +Jڽ&MI�u����?�o��t�t�WI6�	|藳��-/��cXy��]0�-�� I��=�SW0G��SZ������[������J)(bAfa�,��j�o�Fڱyuw�d;p�-|5�5S-b�J���^A�-OV;,�d��x]W֟i��O������G�$�Um��po�������B�bm��X�Jx#z��1 ��O
��ϫCMf�zn�-���"�BX)�KA�wr4`���E�(�� 9�ZmqI��.]H8����7���F��:�� BT�
�=;�ɜ�C�THB�P�����+��h�w�"䐤2�US��U�wAm��;���� �-�+�O2~�V2)������33��S�?\�)0�b�t�1�HRq�2~v�l0���e3�? '�5��"ķ&���Ojh��{��?�a�s{�d���K:w#Cϸ1�P�<�	���GgG/2���5��v*~����nr�c��N�|Nh�wPT�iz��-y:���n|�NB�ڭ��ճ��u���J�c����'.+DK���I�_������_�*�pt��U�e�R����H��O�#=8�@�4;�y�!�\�&�n1cɨ1�㱘-c�X(k�$��Q@0�M���k�O{�"�̇���X�y����=2��Z�.zFly[���@ԩ@��#�B��ͭ�끪�vr�Ł��:�k	#��Q�gJc�P��m��b*�Xp�e�)^sR��]1�1�4�-̝t�2�����zE���B=�����{?vW�TFc p��Eţ���R�i�bX��-����|��F�#Wʱ#hl'}GÁ��hg����N8D��[���o��o����������%����рǩśj~tV��Ʃ�{1`n�0>��K���К��Z�U��ꙵ:3i^�i��u��UUz�BɄ�����AT��Ā�����)}T*�yx����ġ�]	u��>���
�����2\���%�E�4�i%�y՛1SICQ������h���]T����Q�%|<�y+��mU�G�Ҝp���v����V{D�Ș;�QT�-���?�U��b��(���"����b�B��Z���p��~�����?CU�ރB��!̕=C+�oX8��h�=5��2��Oa��;W�-�%�6H�i��3��˔�8k��҇۱�,��a�7-��s�	�:�B� ﬈��H�{9����]'a������7��pZ�lO���b��l͔�w[aݦp�mH��Ʌ�� �!��b��ьz�
���s�/���x2��SWF�C�n:�5��(>+��qm�D�x;��]��<Β�.��|4��3�h�Bޟ�r��%J۳B���mQk�f�,T���E�B&���&c�l��,a8������os�kb��Rۮ��.6���v����^��s�]j�"�SG����Dķ�$��기��N�:_]{ʕ^�DI�\��K�nYW��Y�+����#l�G�'�;�DQ��~���א�����=r��nD�"��,��Lbh�_C���㴬h�������J������	O������yNF2៉�����Qа�OX�R�=\[��O�_�(ށC|�+�,aa06k�m�y���+f����c������c�����}Z�<9��7+��=�q'����/
YJ���&b��jGҳ�(D\XM�Fa#��A7��g�л� ��R"`�C����$\��y-:3���!�S�ж.������U"�h�(ш�P#QXZ�"� �)��Fbl�w �^�_7VCL��vS|җ�C'w�92B.P�y��0�uq"	iH%I2�����uL~�+F�:q}(�NSW��xj���>TS�M��U�����+�f$�@�����\��_�:��L���θ�~S}�YWd��*��
*�����Ҧ�:�a`(�TIz�5N�\�~����H�|8E������������D?����i��',Lw�����>�p	 Ŋ�8
5�8���(��+����Ϣ�n��}Y͌NV��?��T�L���;J�5�@!�u$T�e�hEz���(������:�.�aXmZ�g�7X8}B���͠�x{��|[��r�7dRŷ�Н�~`��c9gZ��3��$$�["w3�=��M	�}�sU������_���7�w�уNk���:�i����M�Ģ��i�R�O��������>�O��7eGu&���]i$������8�m<Y���g\����%N�*3�"�XHp@*!ۿ�|jz,r?P�,Y����Se4St��g �<"��+�݉G*�?����"9���PD
v"��c�Q�~�Y4Sw������zdR���%���[>�"���� 5�C� *���N}���-�#��P��
F8�#��f����6�t?m�2E�� ���r�nl ����݅���� �>:�'���W$�\B`+G,௿F����;-@\�֘��Q��¾x_�� �>��x� �YNJB0.�^/�H#]��}~�>@tR5�SP�/�G~�r�� �ի��J�GF�^Ia�U)��~C>d��h�W��C2�Z�ɭ�C�װ���qL�n��+c9$,�jn6�D�hN��:a#p�n[
Ii��h\?�T,iZ�
�_�X#���$^^�����%Vv-H?[������L��<Zw��Hm���1���2y~���(�a�⨿�{i|����Ůr*��j�Fs����3�7n���OHQ
�	Q��Nk