��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��l�����f�J�éy7�=7?�w�e���˦��X��(|�EN��:D�*��{-� {���hEې�_�p�P�Fॹ(����ұq���[�A�

��я��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0�����>���������co�����c���3HrG��atU��?cɅ�T=Fy�[�'����փ�?!�[��B�/��R�\ڂ9?!��-��N��$�j,���>	FjN�O�$�i������tDn[ŭ}����jΊ�)ڊ\ͺ�MO�W(�J�� ��tU���y��d.(z��5�ҁ�[<�T-E�E�@Wt/�ޝ�'�bKU:����t�Eġ�dZD��ygG�aY����x�1��>�~��܍o_(�"�=�L�����NDB����Ϭ���wS��1^��AnG��+�o�$�����9Nj�'ϤvR��� ��A���q�QZ��iY'��D6��h���9���#�1��R��s\�pW����n��'uq�Sm&D[�ӯƬs3�K���(tL�����^�����UFd,+�F><�`����ھ:>�Ø�&8��0�n���d�d E����q�`�c��h�7h��1<��0����ڭ ���E0Cͦ�k+������e���P�Vݣfk�T��R.gJ�yq�A�"����v>��;��<��5�5��|p_1�j�_/�,���A�����ke�d�Ex,s�Y�q$tL�F���~1_h�H0�����fٳv�70����T��?@����Ѐ����_U'D��BFvY�ۧx�9�[�VM�����M׽y>`7ď�p�O#<1tp���b.���O�"�7�ܖ�[����װDΡJf�72fL�k^���W�B���G��ˁ��~q�ɶR3(�#4�����86ؑ��;%�g�J9FDÕ���Vy�5?-y�}
T�+#���J�8��\s�P�����v�U�j��h�p�Y�������꠿����A
�Q�Y�og7���c����q�,��FYg�IO^�GS�͘q�d8=e�/!v��b ��;���)W,��i��q� �P%v����{D�͞L�&�'?'����I�D��}��DJ�H�/����tQ2_������P.�P�����ΣT�-����T��6z"���x�P ����8IKFW+�ӷ-��)C�mh�ѿ�*?b�x4�"hB%x;D{'��
���@rq(W���t���������]���$���^���rJ}u�]��;��{�s�*9y��ڷ���t��� #!��i��"W��!@�7N}�H���'��d �##��ѽ���Z�D�k���T�rT�7���1�[�ن�g�����-{�.�M�J9��tQ�M� �ξ��D�gbP���4�#��w]���c��%M��[��eP�5�����+C�P��_�)�Ԕ$u��N��'!���p�'+p�n�"�)����a�]q�~% ".�'`���g�Tޢ�H_�9�ʃ�������1�g��=��N 9�,�����D�+�3����2�i���Slβ�.�qd�B}">��1NT��Y���5�?�m�Rl��1�%��m�~�%��5��h�Πx��f5G�����k?���������JHs����7�.��ڈ��iB���HQ��`!?�4Ld��3��pgq^��R|tg	��36#n�������R)�i��P�}�� �{�bPN�*%�ü�1��ڠ5�c��m��6T�|lI���%��'<���.[
�|�ɝK�Z��!V{�ָ�ȲH��puBi��r��(���I���Y����U��V�ɕ�u�)��x�?CS�[2ѧ�ߚp��$�]ӫ
h��?�Z]�^VH ��{!��;���]�{�6�j���=t�$�ЊC�-!_kJU�I"�*�8�jl�������N�cMF�t��ɒS��xv�s�~�o���kuy]q�;a�BL�ڗ������Jo���v�<�Y�=��Jj��	\*h��П�#N�*�b�V߭�},�k}���TZp��y�A�t�o���IpK��;R�������[�=�����/�)�'~������$�d�C���B��`&�}G�u�y��E;p�?Sگ�p�;b�@��Kn|!Ǒ��޽�}�����[�LO-	�<I�Zl4xt�<�U����1�����>���j���(P?�|-�V�Q����B,_�����آ�#]]�>՚Ʋ��кD��B,�N�5���I!�Y�X��@�Ѭ�x�����㷘��R�����C��ю�U$6�"n��. �C1�`�C�X��PA<�%}�>ޣ�����-�K��j�F9����A^�dl�pGy7Z��łs��$'EII�@�q�\�p���w�þW�۳vt�<���kD <��[����(�r�ǚ��8=� ]0�J�{�����i�B��NYX"\�gĉ��$v�R)Tu��7)>�&y�����D���<iS�
���Af?�]qÞ��r2B�18i�UX��z�MYo;���2x�:���{m4��XC�Y�ULC�
�p�c^35��D�y)��'���|V���bqhi(v�?��y��f���Q�y� �G[�:�PF�/�	Oo�W/����10�0��lT�
rvı;'�����K��Ʉ[�h��v���cԗwF�Fm��Q��KM�٬�{]���>s�3ɭ�9��9�����:�x��������q��J|ii!��^����z������=~�����u����k>2���u�C��S�ߵy��Ĥ�9�f�iXgs�o��6h��f(,[��Hz��lM�Ju}���5��I�躔b� �f,?�A��UM"�Ѯ��i�AϳY��{g�p����ɰ�Td�Y?�9�5�Z�#6�{��☴rP>">����>��7i� P �^v�����T6.���9�:�R�w�*�+b�w��0����� �N0ѕ��?9��\drׂw�Uk���f����L�OĜ�'^":��h����ꈓ����IVVJ��y�V+��(��d��G����С���=�WK�i�̓�c����XO�S��=��nS��DU3>լW'p�_����Y~��{P�
Mx$�ɧ�J���������x�u�tBlQh��Q4���0�Y��� ˱
����HZ5$��T��p�K-��|�2yPJ�O��70Ն�����w���6z��q��V<�I�/�뚟����"�m���Q�BU���$�0n��7��#=�ڜ��_�$T	\�hF:�#��]��Y�O�8�O���F�,���ص ��P�%s�O�nL	�V�\/rM)�-��4��X�M�7��%e[��bl��Fj�u��(a��d�lN?��a3_�G�:�$��I�cV�V�aC��.bʹNu�xpYX�@�C�I� aW�f蘨f��R�o�+e�ʃ�����<s��4����;�Q��-I�,c����ΰ��ߙÔ=W;r!4ϻ����?#�ZX3�� ��(�J.����8�q��]㯥>���lX�\�"Ѝ �\ᾨ���u���"�v$�������Vg%n��%ݧ�K�+t���ʸ�ʩFrJ�pJ&5"v	Z�w��ιږ������$k�vG\]bY�%t3w���G"P;�=<�9��Ю3��V����R��5��y}X#]vK��b���u�>��KzZŻ���pP����.�u��������@W[B�zԀ���1�_�����Z�)���V��z[�&Ðر�C,sl�$������ ��偽�7��7���|\��O���h��{�;����+�NCȢu_�dӇ�]+��g/�w���!�D?�6��Q�~U��N���<ŗ��_�K�)��4u�����a��d��S*�§����f"��
���}"�L����4������k�~wc�m�BoP�2��e���J|ģ'P?�3s�U����<U��"��M�7��j����u�~�y�S��3��/�SѼé�֧Ex	v	1�~2��ive�mڛ�3���g�`��8p�����U	���=y����K�WȞ��'�vp3����]8�V������7�_��yr���e����1�X^;VX�N����b?%2Y��Ħ(��2�@�U`�=���M�1@P~��#zR�x#�:ڰw��)�1Y��haA3���/J!Z��r�q��,��;n]Ǐ�%���F]XPnR
	͐�F�S��:��>���s�I?X���3Eԝ���N�#JLY�����h��bE��.`��-�$k�|>T���8L'����u�2����
��LQɍ�a*N����)�����Q~n��ԋ~A-K���K9�Ѻ�Q��D�����[N�@��c�m��ݰE���u�0��/��v�0B~K�p�����:}�Exմ��P>��e���(��l�3�������N|4�-_�F���M@RD3J]���wBE.�i1���D�᪞q�ٸ��	�ѳ�V��,����Q`��Lꚸ<^�jR���>���mM<�#|.��v��o<+�Ӟ9��e�K�����d�qo�ⲍ�_a9�E2�u�"��:������!Q�hgROpy��5��wS��	�lkE�LL �)��ld�P����\��N�����&�K�j���1&C��\tN��h�a�	���M�s�틚�s�(�wpK�a�g31���#��i���;2��*_�R�|B$��)�����?0��b�c@�X]�2�>�y"�J'�p-MX45�v���	6�b���0���=)�e����t<֮����|��vLqg�� +4�K؇�G�������V{)�&�~��!�����CD�&�R�Z!4FG�
�n�O�u���[a��r��dG2�/�}�V��� ����Wy�eU���R.:[=�z�5���W���p��
�}��!jO`�W����<�I+>h�ti�����z�Ŵ�i�W�jf��@�>WN��/�kϝ���+�h#��� tΘ��C���Y8��$2���4PCb����L{B��u
MԽ�m1�8���2�D|$wM�,^C�W?�ң9Iҵ�{B�mP��'X_�A5���y|�,9VZ�VOQ��H�ũ9Y������`8��r�Qߪ��;�>aU)�ނ)F�p�����>��j�AZx�v�Hs>n^	FS�+�����G�	�ì�vrN&.�=	��<nTξ�o1�ե����I$R�C��]!ȍU���;ߝ�A�Sba���F���pO�䩊��ht�x�"󈭜�������zvn��_Შe�~&�ۺ}����a�`��A.��4vSB�=���N�>d�N%d��Ovݍ#aR�0��_��Jz���?�om�������:s$p���qgE�M��
/�$�%��1�М�5@��A���Qr
�=W�E|��旅̀��^��1ڴ'���I���2�~�煃���g�^�� ��0�>X��ݜ�[W��`x��T7
`0,-�m��-+�`�lOϮm�&�lϐ�'�Q�D�H1��*�ߥ�&�����UCY���J�<�
ሂ�*.��~���K
*��Yp�М�I_���U d9���8�
��R2w����6�8����9�V)Â�:�e�����A��V���M�h����8�Z�n�MRE΍�l�8&�;l�f̃H�~��Ŕ3���K��Q�_�Y����Έ�bKMt�:wX@r�c����3qb��Ec ��&g���+�tw��;~� 5V���(t�$/n�{5�)#���?4�>_!��UC
�]�z���K�����#�k����o��/M���ڔ��j~�Q��lyr���9��и�s�9��I��K)G@�p�;m����b�'W�C�!��Pq���>mE�F���#�w���I�?�xH�u���-��p��6庩�`�s�,ǰ)㬥f�CN��u<;&
z�A�]�_vț�>2&;��]�Ug�R��w��pA�WN�>(H��d#���O�P8G�$�$H��lj��)\��A��q�l��9��,�7�'�7(�D��3H=�L��%jG� �ե7_�8��t���͇�4$Y'v��J�<J'Қ��2_TW`g��������k�����
�;is"�`u2�����X��CG�u�'��8��y�y�"�E�����rL0b���~�e������;Sk��e�����Yw�cwfz�j^���{Ɩ{b
dW�Ϣ(�Y��&3� ��1o�����,�1QC���a��;���!�5��B?�K�lk���xO>�t��?�4��9|����#ym)�7s����T� |�Cw�.
� {�� �%r�h�&'8x��З��Oն&���c
ኍr���5+��|��׷Rł(���W8�⌸�~����=�y�3P�;�U��ѴK�P�&����QQ<ᱴ�g�X���4\3޼u	Q�@14 ���D�`�ĸ�n�Ɲ0T8��.��.4G�ƷY�YL����˔~��K�A�?"��C7���a��� ���STt��R���$NVɥi��;�0kL8,m�?[�ZZՍ�Q�:���"��Hٚ�M��(�:5����^7�8�M��{�d�!|6~P�'�a��7������]�H��\�+�ϙ��Dl�J�/5+(��
	Խ�*��i���w���u��u¿�q�=
)����;���|��:�J܍H�SqHyS�u\n���� �^�o��T����t�Ʌ۾�}���}PE��feK� '�~򵹐���X��"l����1 CD��^���A��Y��b��c��o�B?��ko����N�WOǝQ�Q�1��8o����꛶��f�K"m��k��C?�zu����:9����D<	k馨�7M���:�>�L��7��L��݉�K�ފ�&��3|���6��\�`�8Eg��(v��v��M�#u�63d硳:%����['��P]�έ��Fn���L��+C!d��B��-'��Ř�t��꫺��H��9�e�[z����	�N�3���_*ԲR�˕�d˪����x��_x6\��=��wͬ(D�jx�?M���+���ma���>��˶Zk�BTB1fm�l��+�����C?\5reKw������]�V~�)S�~�	���}Ȯ����oΆ��E�d*Z�^���Ka#�X�''��w@��T���ؾX�#������s�ċ�O��"Cw|�r�i��$[��n7��]e"��j�_Yл���S9V���p؎FPY���AEZ����bx��0�ѕ��3C�U["}�bm���=�X�+N ����3��д<�U�;}f|��q����.�����-�~#R��d��B{����/N���'�
Uwro3�1�2��U�[Q�����C�T�K<�KE3�O��?�f�u
z�ίG.�����AX3.�@NXC-|k���ٓ���M����
oP��l	�E��5N��"ᨀ\�ҽ`���t, �y�A����M���1VQQ�������(����2�-zdɕe'�J�9��J�4�B>o*8� ��R �*u�G����Z[Gb2��'�J�����W�w�Ar��/p$�Q��D�k��lNq+�Z]��
C�;/��jI� rj��kl	b8X��ľ���1�%3�1��Af���9< 
��=L/������8��)�b��u��|�s;���X���� ��`�%|ac�#�m�B:W�b�B/W�=�]g���d�eYx\�U[s=lN��v���/)3Z}���
�
I�	�x�vJ�}�Bk=��x����+���ā<�J3�-�;~�Ϩf� 6�	?��ɞǣ7��J�H���m�>���y���4�ya�]���7��	��~�fp���
�-��n ��y1-�2Y�����Ɵ��(T���ݜ<�o��=U�-m#9'��%�ۼ^�t��;�^���Xi��:B�#���v>��%c�JP��2�����P�G�1'{��IQy�:���c_e�(+�
����u�>Q��f_��B�>>�E�dg�0���j����n7�٣�8�'/�\����j]�Y��������.��~(*D��<�	�2�P�Z�A#%�LF6#��$PH{�[n�0��/D�i�W��L�����;���r=0��[җ��h0�ʚ�&�&�Vo�а+A�$u6䗐� �p������̦��w�9��@Jl\�G�����#0�mtʔ��T�</ـ1�$`~��;N�r֐0ܩD���K�p�<�;!������􊂇�aCi#�Uv}#Qo�J�)^�GNȬ�+�%��4?�v�T�ĺ�t��]x��~g��ț9�Hx�����a�f���d3d�v�_BU�f�D'�f�/|�Uz��B�'�@�����ջ~���$��b~/�i�He��[��O3��z����8	���2o�W?����(K�F6�ۀ|q�io�0�Wж]����mG��������ʅKSڌ'���L�b�����yI��-�MH��"��O�Ґ:��2pj�����O�����O�X�}wd�N�����Y,���9,� ݐs{�6OD��R�.��h�$�'�-34�����gಛ�(����A(��hv�3����.�33�Yʯ��:�<�2�&ѽF#�qf�q.�_��ϑ45inܘ�GL��1�A+�
AW�PT& |��ࡖK�O�� K����'��x7K�vV��U�
Z~g�@�N�����f��8�/��믂���1Ӫ#�C@'|D���u�i󑲉0o�S��n�u{ƙ�;��+E��|�|b^����"�h\ν�P�W�IG���(���{�-��JZ
�X��c#��aފ?W���c��4V
9$��fF ��F�%�,�j�Fp��Y�c�
��#~��ou%�+�}n�롬#�v_u��ψ�\ UX���EV�̀q�>�0�[����Ӣ�	ؖX��[$S���)��H>\���k:��$�����u��z>��69�f�0"�������ૐ�?QqzDZ�Q�\umc�ݰ9l}8|]<�!��N�g檱����F�ώj��G�\�����޸t���o�.�L'FL��g�̼�s�>[�-�Kh5>h���wK"��g<����z�Y��2(����|��X� 
��/���G��fߦ�m��Ǯۇ
����	9w"P~�L���͙)(!�5Ē�Y�Q�b��t#� �G�8u���m�UH�'I���͙0El�دI��{[�Vx��K�?��÷��}=i�P��	:<7&��<}��%x�r<t5�jQo���,� z>��M%�i�p�$�81;2
���4�ϵ�2�p-w���<^�~���x?a0D�`�����J�����rdt�Vё��nЊ�X���4i{$��b�¤�Y��f��Y�+,�!f�� r��(�l���1�
v��s�z����÷�����Q�R{n���{�3�a8!�Q�D��n�i�9���W����Gqw�6&6'.����?Wq�5й2K�@�;�oi3ֲ�6jp?�|��*��5�(���i0B�Eg`��� Bz�jg[=����c�!=�k.> 4�酒�m������8?��f͊6 ��ꤟ�eխ'��OѹV�\�r��l�ȷ��6�&���ꝃ*V���'�fT�L\�>�L��/�k��ڒ�f�nJ477ۆ9�>�Wi�aR�g�C�����<��(��]�����Bm˒4e���ێ��ޤL������P�un� �ITRs/�w  x���{�^$�f؛��w�ɠ��ӧ�Ʊ�z�Qӡ<��LLI|���0�����H.1��Yd۲aJU
9���EwW[�ض���P���X���KԢ'oL1�hԯ���z��Vlq�A��}�5�E¨�7�=3p��Xߠ��WP��J�SM�EwM�T�/�t�&�Μ��1Q�X�Tw.>�3N�:��6Q+����b9
�ç��'ǯIya]�r�sHqW!1�� -_��G��A���LZ������\:w�D�w����~GF#SF����l�l�{bD���;?]8l��O�_�WB���_烅��&��%T�����0�����Z���v��|��-�����|ϓ����Oc�#�p+��751��Ќ[��:Ӷ��Vj�ɛh҈�N�	�$�ÉϜ���k,��'>W��&���.5&]�­MD�<��ZԘl���/�j!�BݕB�M׀.�P�.��bC$��a~�&��s�,�z$b��|&	�'����af�+h���!���w����\����y�:�žt�Is��W�����&K�:j
-5��K�@�$N�m0hx�M�EQ)�ߵ��lq0^��aT�J�3�:1�4l���M�u
���y ^71&	��pu��=ܪ^�������{)�^wX]:��U�V�d�:?eG�'��y:|eR#�������/R�z��@V�*#��Tx���,�>��Պ>7�4���������j�OTE#k�SN6�n�F8Ѣ[�I���'y����3o���?��㎦Ӣz���FX'�܂�E�y��$��������tq�g,-e���o�T?"����Ї�oi2Dx�z�%+,%1��O6�o9�vxz�ʦ_U��Υ^^q@�;x1T��R�
���ؓ$�g]�S&�~u1�hUf���~ϸ�Ѿ�\�O7�bɤ���=U��@I�&_8Q��1~A��g�\�_�)�fř���|>!j�[y�20����4B*�c#�/�H��"���SO`1�8ރ�.:7	R�.'��������B@�e}��)��w���KNz��?N��w�_�3��>3�xsM�`s����$��VB��z���6]F�)gx�E��ߡ����&��hq4k���C��Z,��ɚpD�5¡�%:��78�G�ւ!IB�@�'�X���mЈ #��;� O,��3V�Eow:������O"���s	</D��aZ��M���T�W@������1��k/_��%�������k�'��g��ڟ�v��������t'�[#Y����ܶڎ�OA"������0gB�r�R��w���c�J8��B��Y����7E���
6(������j�߭�
g��ں�8CX��M�0X��3\�#�"b�m��cp[�F5�`Э��Y����EdU���{FM;W�ά���ϋuj���sKy�v�Р����iĈ���ͅĢL9n(��w���􂀊��w%��͸cC�����g�Y-p`���oy� @��nI�M� ��t�����m5�񯙃��M��ħv��Bx�VvR�F�C`-��{��
�<T��"4q�O�}��☜��d����-�F8�QI�%�z�G�xIj���v��[��
�zLth��#yU~��T�A[���7�h�!�%2�*g����B��z�{LhOm��_26��o��{h[d<�W�YC��|�|��\b)��Ai���o��я�
�m��^"o0�
\�P?����)f�X,��$P���bW�ʷT��g�/◻"a����Xr�/�\��t��I�mŎB�"_I�z���1�;�O������<�����f"���Ҟi����Nѵ���RkK	�]q�q�xv}�1ڐ�����k�'�c��>eT
��t�Τ�l��m���Yg��C�����y������0Q˹�T�"vGi<G�1 �S=p����6-C��̮l��!��r��>M�Ek�,V�F�u�L���/�.R�=�_��f��Go�pqB���"��cOPY�u��^W�G{����,i����$�dEπq�N��	�-��(B�P13{HD��s�����u��vX�&�i���8��s��us�AN$��6�,����+����ȼ"r�"����Æ��h���^�2�i=~���P�uBs�?�S���ؘ����l��]�G!;��A�ࠝȉ>�8+ˊ�y�zNc�y�S�c�H��p��A�ug�?�a���ͫ�M����5�*!�����R�!��gC��s9T��T �Fl����������O\rne�x�t�Eą�$�W��Y�X�W:��W�Ӽ�[	���0�O%���Z�p>s��6uҟR^AQdR����4ǵXٮ���<*E��@AۂTj�b�ݒ��5�J@�X���S��a���'I�,�p�Rd�x|)���=:��sm+�vR1��v]cޤ��#4�&�ҍ���l���"1�0n�"?��(��c�����	9���[�+.Z����s$a'p��ME�Ubx4������O4����{ �6�9
����mo |�Kgf���vb�[&����22#�~+o�۩���QH�����0_�Byαo�om�
���Ȳ͂�c�)��տ��O>�)����I�z�Z?�s����&��4ȁ&�U�|}Y@���WG�4w��5Z�C{��A���� ��|��|Ay(x�;1\�h;L��g�a���%zN� ,���NV��h��z5���<��حZ��!t�ֹ�Ef�m�h&f���A`��'D���`ܖJB�	Ǉa�l~���
�Qjj�� 4p�Re}����j��B�"���T��7k3�
5�[7P ��Hu.(��8X/R��H�X���IZ�F"��Cy��8�m(���0'.5@�����L���̍PO��N��aW�F�M4@m��-'�ζ�Ò}k�]���"��*���738ߋ�ӯ�n6L&N5�<2
xh�Q�:f���a3���-B{�{0겙.�ki:h���a~��ڱMfe��_ABAI�1f9�-����I������eg����;���;0j092�Sǹ��x�/���d��>7��CO6M���V-�C�[����u���p��d&��Ϯ����:�|5Mɒ��d�Ԧф��6 �b�Zq�l��]`��e ��sB�j�K�Q z	���i����_ڢ ���]ȗi�ߤ��1�>�TR����Q٥c?�R�H�F[sW�=m���E$R�>"0����x�#Q�#K'��%/�O��I}�\�\��'��"Up��D����W{��E�/Q�嗜�����=G�����#B)K�:�� ݫ$��rN�C�W�)&D�`��,��<J�/������k �����kx��,����ꉊ�t�f�.�z�D�?*eˋ,��_�n�iX�R�d4f�j޽���uXM!��ň͞B���a>!����Xf�Whs\��FX,R+W���ۣ����Z��fΔ@_Y�j�tٯ[��N�-3�����.�*����0Z�|�Ŷ�n����¾��g��e�t./�[�|��T�:&�#I���3���Yස�֨X3Z��aU�?� d����U��@�c��M�;*����m���p6����Í���OaJ�����"A{�AJ�-�^�IP�!��1��̯E� r4�i�c|���Ɇ�^	��L
kd2P[zc,,��㺽\�p�q&�Ȋ�=Pȏe?C]=E��?��㌉Oob�`���ڥ�h�Y�6��-/Wf���}^I����W��+��$�؁��$�qҐj�-�����K�jL��+����=RcY�A��U�׸����Ț���t'^��|�ǛTu3�0y������,����clH,�q��`�e�,.[�54�7��W N�����4�����(B�G�����U���K1��A���J���)~��p�WC�Xt<:	�&g�m �4�v[Z)���{�j |E�0�eЁmx��5о[Ӵ�	����������t�{(ؗ��4x��"����A^��:Km[c��o ;C�cNy")�i�r���8��M}��v\���
��
I�C��]0����:�O_�<1\+t�,N 0�6�*Ί�^��ν�^��Rs8-��% #��M�A�>���K[���˵ĩ0��gn!8��voͼ�.��b�|v}>�3 *<�%���3���X��nE� a8��2�~{JM��x�̬>�I����˷����k#)�/�Im�}�ߗe�}�.o����;H�v����^��bͫ�خ����F�����O/�y�����U@G�	�)-ipn,�� Q���aze���i4���m�8�i�K��c�Ұ��W�ΎHjJ^����ȯ�IB��_�C��X�"G�i�0�����R*1 ��6�����K� ]�k��ť?��h}����½�f3����h�V��X����{{��'���S��̃�0��,����ff�{}J�v"�i�!͇�?�~��T�%�Tps�W��PL&�i�����5;�DO'�*qw���_T���G�W~�
m3��L(�	K�7�����Ox��oK	!��u��C7-=�.��Y���858�-�0C��Me�6�ˮb�:D�`mj{e������/;�
����:v��%L_FW�b��ETQ�s�(�@�]a�,�ER:PMu�z�ZAv̄6Y@��#�m��Y'\9SQ(���	���j�G�����ΥdX���ꞃe�`�n��P9�1�|1�����λu�e ��8�g9M8����.�� ��,W⠧:�V�r	���f� �G3P_[�k��r�N����ob.��E�	��(%���i*6b�1� ͯwqFQ�.�aΦg���-	���#i,����8jm(p�*����%I
L�l���'����D�ms�٪sd8uH�#�)�4bԙf<�lދJ �fO
8���k�rH=��Feӓ{���n)����N�M����c��I�̟ym@�����J�dQ������O# ��^�����Tq+AP��S�']��%�%X�qv�
�X�`SNb�Gi]X�g���K�kϑ������a���'�a��D�Bl�4�TiU�m5��"�(�\���KYا݂����-<-@��-+�>	eNn4ʖ��G�[���ю;wM�a���( Y��!���ϕ8'?��z�����fZg�5�m�(~�6�Cj|:L"w�1,�#}<6��#]��eWp�;���,&q�����%��$�זU��>�������6|/��~A9�������ȏ�cn}�]���TG�.�p�x�*�{������EP�-F�gU�m��[��h%w;옓���K@��!M����$��UU�����-
۫̨W?!���S����� ��@s�X�gj+�SZ
.v!6�`����>�K���SYj���]�s�w�����$uo��u��J�fmmjU�y׽�IUb��Ғ��$ ����������_�N��T�B!c����Z��X�u޻�~�N���̩x�FSP���o�(�)�<�E�p�"���K�w�^��AJ	,&�%|ֹS�
�g	Dxt��+���7)J��6'~7n��7��d����.g�u57�\�gKV�3��~�����O/�U�8��$�k00�npY�e	"�K�����N��-� n�-���pbM|���f.
Æ�6�[t�M���N��|Q2�.F`�S�*0�A�Ջ�VD= /��2ص���LNEw��fT*w��J����a�glb�(�{�$*��H:.��}�,Oc�^D3�R��H�n�%Nf��Ɗ�
se�F���R˘��G� ��=�G�����q��N��~�F��g*(R`{�Q��_1s��q�ԒOehJ	E�y����ϼڏKk�F��cf�����]�|���L���zA��~6�]��e���uT����jM��:@z` c4Q���a86+H����9u��5ut\��|XSl'����e������
��v�0������d�%�֏�v�Z�����<�J��E���Fٟ���$ ��C�Z:��2c�hq�"ۛE~�V|'�1���DP2Y~ȷ�����П�EK��ף]Z�ƨP���c EVf��)rp����h62�\�}##!1�]6L��ѳB�SQ粖pܧ?�}gիr=i%J����l���;y���-B��;2ɜ�QSc
���D����@���Ⱦ�>�8�ӡ aL%�֛ئq�Р�s_ V��i �%�I$@ek3���n���+���Uf���쎭��6�t�To
�0`�I�'4��u�ĤQ��>L�ts5�C�-!h�x�� �`��4ܦ�㘋tb`�6o���!J�ɼ���𻘈7K�D��2j���x�D��³�޻( b�Tp�!^2��蔢��-��ay�C�����k����B,�����9B���~4���8��� ��R��H*���1�M*S�l��#���kҙX �خMO� ��fvY���.��̨_��q��1oXq �|<�2����v�3��UH}==�`� �����G�!N��V���p	���"����M���E�ULi�@���=�MgR	���W��+�<+y��Z�� ̢�c���� FSAmu�u�0rG��X�4ɸ�7䶶�B�-;;K5�$ʭ�@:�{�j��t-�pЬ�ܕ`���T$��3�&��ia3�.vP�O,)S��}�΃��B���BSA�ĕ�#���U��=�/D�mb�����"�J��]N`�2kʼ�������%��)cg�-�|�&�iS����UT���^4��,�n۾�p��(i���)[¹�hUzDi���}��P�gƕ�O�I)$^y8�L�i��_�1��8��@�_6�۰�]��^�]�B�(�!D��
u�,1 {ٙ�(���`����w�r���(��UL��-�aM?�ĉJ"��
����v���^ȴ��`�ΎY4�C�&pZ�#%�k�R��]1���3�ۦ;-F�y�o��q3�mQ�:����[v������4f,Z����z����\����޹�kf���k�j�JM�_���\��0�I&N�O�n�7󯣐��Mߌj^9LT@��Q�����Ȥ��X��T}B�3����`��{��`Y��C��|� O�	T��BO��V����`����/-(��U�r�}������P�� c]���Tީsm�e�x���)���4��r��XNR?�d}�S	N��i�+�TZ0iRH���I�ih֦c����{��܀��A�`��{r��i��	S:��'�nFAq�A���F��D�$�^0^ƥ)��JDqeu�OF$5��(@q�ܮ�L~��s��I�m�`�Qn��i�+6
��([�Ѿ.R�税��t)��&�S�CW0�R�����:"�o�	(���E�{��U������|�Uƫ  \�:�$� 5�{��υe2�t��D��$�3-G�$�@�O M�^h[{��U���o�����b��ɵ�-��:���t:��ޯ��?p�g#����W\����ґC54K�@�Q3
�ݺ�	�vx��^&ӛ�K>�2�Ƴ�+3�h�sk�;Q�{��{ib|(D
e�K7�0�;m��Q�����UF���*I_��ǝ�=��H( ,�-=s��v�����@a�J:�p��� �dL�<�����|6F�^2�#�lE$P��J�S��z�U�h�Cz<0i�gc�lз��H�g�L�dç~�K�M%�,�E{�cx�����(�:̸�I5�����%�β�$���͡$�]��*yX�+��	�J�����
��te�"�M�:u��9����P�;�����Yk�K���M̷����4�3���F5���j��!�B��O�ȟS�a4�yr���0)��cw�i���ݵ�ۋ�t�M`NxR�W���@S�㖎���<�e��dD��M{�M_�]�?��}D׮��jۓI�Y�@�`uSy������� Lv��7y����ǧ�:'���֙4������*	Ӵ���'����{;��Z�ϲ?����~@�V,;�݇\��%�L�����v"�*�Z-�x$�R�05Q�� D=�͵W	�~)U�89�Ƭ\�)���o3>�<�ٽHk��f����-����x����7�F#$�d�{V]-���.�hi(L�4B�(�v�8`�a,�EAHevs07VH~@����o�j����7�o����7]�Qf��޳�7�/�K1��Sі$�D���>���9�*�yg�BOP�$=  ����R��eա(L�~	�X�"^>��q�n�UM��8*ʴ�s�������T��h������:��_f���8d����BD�����	�ڨ�/�@
��$,hY��t�e�5ʺ=�)�L�u�*, ��PJ�	�AÆ��'�Һ$�i.�mk_b���j���i�ЈΌ��3���<��Ҭ3Z�p��?�����OD�<|y�[��2_�ƣ���4�^��ڌװf����s�D�P��!!�v_��~�E*L���u闏�c�W�y�3
f1��4�������x�������7K+y�ʏ��ݑ״UQ޺?��"�9rw`�^�$v�!�)�SWN^�y~�
6�Kңh���'�{	z���3tw�9۲;�Ah��q�kR�ޟL$��\~TX�h��%�I6̨0Xof��J�o�1��P����v&%�f~9ˇG�i5s�Z���"4�tF���(�6�rv��L)�9��Z�|�՘�F�4E��d��}a�s�������59��3����&u��Ͻ$ʶ���c����h�bl�)�e��0��I��:C:����R��\�N��1E�/�q����(~��x?{=h���m/��9���
+���s`;y\y�l��@4��E�`�G� �@8�^�����yX�>��PY*�z/���K�H�dZ�UҞ��]�:z��?��������]�N�5����@8�b��E���Ӳ�R���-G��b} D�T�.a��%����emBYb]?Xf����tX��Ϻl�����)��^vJ�}�[�LI�0�H���^7e1ް�k�/m�4��k��x�f�Sv���w��R��au�T��A&�W�˟76�U$�|�n��xp�Pli�к�8�p�ة�e�?X�"٢�ہ�[��a�x ��Vx�?����i��'�4�4|�!s���XCq�QO�%����0 �Ǌ|����KHe�^��\�4�f0�
R�y��n�lr�
�PJ���F
���r8�~�*U�֭,�!��=�QѪ`�4DUR����#�w�-.1���/y�.+Ga�7k����pۚp�W);Ԡ@����T�fQp0�t��d�W���$w���AǠ,���p���h�de�^�
�s���C�G�&I=��eP�X$�:�n�n딽L�}D�aKdU�N���>�\8�]��F4���EY3
�m��_��e��J�f{�)Á* 2i6�Ss��d%�E�@��2��
��u<o*�˻@ݏR�1.�/I|P�`�D`!�U_<��p���K4������e&�q�Z��$\z�g���-�k��:�8����I3D�R���vBAx'��@�Y�W����{��@�����Y��V��G�&&�+ ��&����t�v��^,��KrO���1qE]����S��K�}�JF�V�/t�N�$�̦*�ؖ�r���$KE���*x�z���KARJʓ�t�' �L��ii ����P�sT���Yo�m�#�To9A��U���X*D��Z���/ƹ;�GLZ����/�n�!"|�G���~�S����������}U�i�f�Ï)����z���
�f2�~V�����ѕ���Pf��W;��,�c�G7`�����ho\��y�m̄><�OɄ�w����7+c	������~J�ܗ�W��RdST�5=H���%7��{t;� �kߜLʃ�>D�V����l����ܭA0���s��1y*#���U���%�4���˳��r�K�ʩ0G�S���0�X^V��*P�D~(((�nܥm�6��~?I�G̲��R�y@"9яx���R1&���90o�����ytY��im#C���P·�)@
S���$@�d�� J�֛�3/&��H�g�J�%�t�
K?z���D�M>���'���������D����>GHTs~����. ��R�]���0�M5ژ��V���IRG�m��3|�
,�1щ�*�U�T���}>�<o<y���&G����c�G<�1<��EJ��^E~P?s��Rz>��A,��Qe�|{X)Q�l1k;ƍ`��>q��7$W�%�$�Nx�<=��-~�eI����+P������l^�P��$ '7:���i��
�~'�_�i�MEz�#���(�*4
��O�K�@A���G�j3�d��z�D��&H���`�a�%a��b�(��&͝ HW�Bn�8����LH-E����j�g������M7�K��()ſ��҄M�kkJ��#GY��������1M�f��v;k�)y�ͩjl�û�%����5V`~��|w ���ʖZz�L�Q$��EJ�XǄO�f]t̂���|Iߢ(�8H(���CyNQ���-���X�J�*��&���Xᯞ$[�F���06�u�~s����tX�`c�B��n��$�V����2|0�q�@44D��-3�E^�}R�BC�����tj��R`���髯%(�R�ll-���t2D*��!t�_Ǡr$���3!(�fJ����.����C��������M�Z�>�^��iB�H��ڞ%/���>]Z�0;~d:h�p�9�y��Q��2���q��`.�������� �?7E��I�ceY�A�f��9����.�ȾT���.j���6��o�_cb��k����̒�����-��6����m�Q�O�"��V����j�C�"��W»�B��vn�l�(�.m�y��p��[�X��S��gO�
��5��d0Z���#�eI�g�*�G:�����{2��n䈚�]}-4�1S���� g�c��\+�jBI��KIi�)o�>A%���#|����f@6&|9�ҥ��\��O�p~atX�O�<-����zi�p�Zl~�J�:WU%������+IC��Jj���`P�?��i�i�xO�[�ĵ��#$���G���g���ŘbF��A2�0��z���HK�-g��rN-�q;8��Z��`q�vY�ߧ@ݜ��+�����J�1ȽΓ��\�eW��I�4�a�zlU�����O�H����
k?�+[��K�F�m�^�{�:��x�G�ǧ��nܣ�@.���$�iMNmd7��"��E)Jm勚�M�i:m��N�{�}EG��l�Cb�@u�Bj�weV�J�F۲�oj��A1�y���P��t�8c��;�3=�Y�2-�����}筣�;�i��Ȇz��:���r�������qI�B�,Gw���Me��K���C���	�.>L�P�n*���;%e^{+=����;8��c��E��V"V`*6A$���@�F�>W&�k�m��W�Ŗ�95Ɯ�����i����E��fn�F���5f���)���+$�i�ǋa��z�����xU�X���Q/Ѣ\�I����<���h����Dq��T�� ��󒕙�}��0v�h�U��Fϲͺ&]q��"n��o8�6lm2qnu���a'Wjr��i�Pf�j��X ��<���j0o��E�O��4�E,�oCβ�7��A|�3ҭX���T��ǉ!���@�T@��mE��hf"W"j=�)T8��r�8�r�����@]�hG �U��R���µgi�v�&{Q�����j�c;6��{��R�(wVE���^)��/�"Ed�L7�!"Ԓ���6�8v-�G1���W��	Y�[`Af���s8P�=�k}���+���!����)��>U�l�wEϨS����qY��Q��,J�E�\�T�c�@��ȍ���������۪f!ITRI�Z�e�����_�q8?�5���s��Wce��z��%=Y��n�=�cZ���t���Q�������1�yƗ���]f�,�8|��j�k�M���~\w�(;�jA^�t�c���V��jA�����a����P���ڙ�r h-״��P��ڡ_V�q�B7�0�Y� ��P���H%��Gf���Q*Z3�f��{���t{&�M�D� MC�� �� 1C..��1~�m���|{��3���D�����J� aZu��˽�b�S����oj����C-���S��;o�,xU޻��5Q���.s�&�l�r�f��^�"^I�:�x�˱[��&[�8ȩ�|���-p��A��4�/������6'�t��@Ic Y��S�+����8��*H�,P�>DN�2�A�#v$��/W�=�Gz꯽z|ϗW�����N�3�O�WSj �#.�p�L���:������|�3A�ꛧ1�pAA�^�٠�JG���85G����0��T�hM��K$M�b�Tw ���3��R΍����f��q��q� ����ݐ��b�jz�+�iEJ��g���`_�ζ�L6������oi��*~p��N/����D��NRt�̬~w�&C�)����`^`<�A�O�6���Fe��E�}~��7�p�
����1α�(���2���
8�ʻG��Z
���Ǧ6��M�DQ��1� �4��4��/�@������M�B
r�a���KU�� �';���=菟�LY��2@�;{Ĵ�D��6]"������!�\#��t��G}~ �~�6;q��ڄ)���Ɵn]x��	�e+�,Q>,(�X:�=g)Jkli��]&[���*L�����q� �����d�.D��a`�r;�$�r�M��P���#�5f_e��`����a�zb �G�������[a}����jj����y�Ӳ��I�q�?�P�l�&UE���� �+	;�����@�),D�2{<�g��V�Ze���}8�)�_n�9{���n��]�7?����"�c�����)�E�o�8Q����,�b>sȨ��$��O~+����Je���L��N6��?�3�b�6��w�xe?������v�W�Nbɱws���	����9 *�pKO��K�z�}�J₵�����V�"XX?�l\f�6�/�c(�7~;��y|S���E����+ΉN^^���.1"�u�c)9���W�i0eGW������Y�L,i�S�_��_��\�ԕz �3��a�U	����7�k&��qxFOV�YD�k�0�8��LD1�K��^�l��^�q̈m;�*�{�w�rvkc�Κ5�V�;�WB�1���.���n�N�
X)�a��<��;Ĭ��1k:�	���њ�(}F/�����CL"8l�"U1��䖁�ށ�.EO��g��:�����U\Ś�����v�TO���C��{�DM������>gƐ���yv�G��,�f�fY�ryB�<m��V��/�扵���ӥ:��ɼm*ș���?� ��i4�����)�l�^TN�.N�Re�6ƫ��A��j^�E��9K��<�J�-e:�n����F� ѝ�L���G��ZaP���ч%���'Gc�wC�6�`�&6F����!��.��Z&xD���E�2X-~��`�r'3�}WXho�fQ�%�Zj+��	����ʊ_��W�Lχ��BPð�� ��V5��g$&!@��-�� �O����H��aF���T�C=8]��<cL��ߧ�E��#,�a�������Z$â���M��xhά��)�E�������$Qj��R��½#�F�~�,eQ!�4Gެ��͜�|U����D�~*�y${u��Q�h-�S�{irʮ$K����Ř	�D��Kt��w1*���Ɋ�Mlq��:���v�8��V,t���#�a{���z(�V�XM�g,�����߾���5�����,��3�2~ [�~�}$��΍�T=%�9�=-�u�$2���֩�;l�(���N�&���px�f�]�-�`��r[��\/5�sϸ%5��&��>*!���P����?Н}lC�9��a}<(�����K�I������,8wyv���4����T�T&j5?��iy��q��?B�>jI�r<������i���/oi�$R�ݳ����O 9�e���DH�
	-�1�1��I_�;h��i4�[��cm��ؙ����Z>b�z�T1�'�Ї'9Ai�/��,/B3��)$�˶u4�gg�jw�x�K�W%�]�ZW����#�?�`�#VkP��P�G,@t��\�CY��A��
�w��4��=K;/�5	�Fc�EP��hpE*����6�7\[��@m\����o%;	_���͜�Q�V3N��Z��o��X���crO!�{Sw���6�=�������af�MT���|�:"ND[����xG�l;��f��B����^5Ӄ���� v�$�h���d�B�X���EĹMO�;��C���FE��Buh�Č�x�Q�%`�~y�a(V�k�:Ϩ��1t�׵�D%�3z�_���g����1y����P�
�.i���yW�-�6�W�+`�Z�+r���:<oC����<n(��!o(��D�ᷴ>�I�N�z��E #�ƭ����@#ɱ�#�A��f�#À���\\�@[�j�qc��P.�1��d��vʀ_��x>be|3_fsp1�Z����1�,��P#s�'`<0	��bǻ<�b���&<�*[��A,�:�U%q�M��ȸy�r�/G1U���<�aƽ���1�\`����`������t5��i Kc!~4�ep�I��ǒ���@ܓ��/L�Ѝ�koV=�ޞ��#98��hw���*µ��X/YQ�_��rk�.@DhZ��_�kI��g��B��w��Z��8�������PT$�T	_sP���N��ã���m�iQw�:����l���6��x)DJH�������ֶ�WkNq"ٺ���yN�BXg=��k�D ��Xz�ݔ�-��o�����f
vn��7ZM]���N>[�K��
5J�k�O�(8�eXO0�ux�*���G�;�� ��K�gE�2�:�&	a �����#��x{�eTq�yk9��?8����c��ǧ��1�<��yX����,�Wm.9��|�a�;`�$�M������_���@M�˭(�&Qγtbc���+b̠�ט��O�������ϥ�,ou�v��
���\i�<�oHf��єb��t���ؑhFi�K��(_�1Skn�B3F�{�a�ɟ�������{ˮ����Pz�O?��fp^��荇u�����Qxr ~��,e���v0դ>�S�r���fۯ?�Q?a{���ӅD\Kb��:��E�e���ǯ��aԅ��c��k7U	N ��u��;���1��t�����Ar!�0.#�t�;E�,v�h�t�j�r��P�)C~N!���z��oX��X���K����`U�H�����٨ef�73��8J�AK'UC��N�-��������K�
Z��|30���:�}Q�i��x�}�81z��ZVn	���|`���LhHz	VrH{]�d�����Ϩ�Nz�yh�'�%�d�4�v`������q���*��C��T;���,U��0�]�����­I�C�vA�v��Q
�t��H[+X���O8���7�a�kB��n���!k��CI�FP������!!�ɣ�-gz��_Ѻ��V4&ǠC���4=>�R�n�]��Z��0��b:F�����#w���t���0m��2�w��0m�ʧ	��Z�P�ZH��~��f�,%��bjxb+�F%����_���q�����_�RmL�FǆN�t1܈�5<�J`opz�0�Quc���a7���.A�YQ&�b�G��� ���,��m�����Ϟ(�&�z�Z)�މ?eZ�|��GӠLi@�:�̊|Y�e,���$=b��l���+H~�iA�r��&)�a�Z�˒`U-p_P�JPr�V�ɓ�pY�/y]�xrD^�U��/VSw)4@[�����ܑ��ɿ6p5�����gb��-���ͨm�>����[���Oi|�����ʱ{�>�w32�|��,S<�KZj��G)*�䵅��CZ��=�?��=�G٩L��rf�~�4w��jV�ҝ@�	��K�1��?-�(�v�K�FJh�V�+-E�1Q���8���n�l�G5���14%�)����uOuk�]�dM��J��Z�l�g���mZf~8O���4��*�z�*�R��$RT���R\O��������O�3��������+ e
9I5mY@2�yN!�{����Җ7`L9��
y\�jT\mT�۫e�@c�Rz�<�����?�Ld�+��]���4�=��A�K��v�Ѧ�?=��{��{q�AF7����2�#hN�e��e��!����~�G�i�t\A��pf��C4�Y��ז��qZ�(�����{Ope��0����7����G\r�Ҝlb,��W��B٨GAq1���|��cO�(q4Pe�WR����LRRR�	9�W+:�sy³���7M#ѻj���[��X?oװ  �@}�o؉��R��Rdc�mw�Ү��%��С�o��9I+�_�i+L��wc�BC,��*�v�ng���Ϋ<�-��'9L��8Dp(6d�6S^�tTw�������!��v�܆7�7k,��hs�W�A��m�9m+��9P����9�)��SU��{\�d�`������l���볘�E�(����?��7~ܵe-"Rܛxt��U:��K/[hs��iR���k����&�����ME�0��@�����\�y��ވ>e��Zw��8��YBNq$�@�!���u1���Ͻg�cIEW�~�iܔb����a�č��%)4��T[್0V,v��;5��������ȇ�.����0��(F{�����Ό�WŢ����`��6�|yO�� j4�\�l�����h��{�Y�7q��
Y7 O?���i#v�V)�{��y�Ԭ����~bY�B�n��ā���w9����t~�d��;��Δ�k���-w�:]�^�~��zwo���V���Y��*��9te��\���*��Rb����Z��	�X�K>�R�鹁�@y����F8�?�A�m��e��!LN�Cؔ��=-"��_���:b3tV�,�3��� ���)P��I�@:\�z����ix�	�^N�K��c<�"�4�Y����M��������Hd�S�.��}�3g�
c�6���|�~���{�6�o�x��h��X��`*�r�-����5S��!s�gF��e�O�1�J�q��VU'�&��nm�_��'u;��D6�;�$�J5�j_`�n�,��\�0PEP���˞�ˈ�ߚO��--��z�5�J��!~���g�qC�*��>�0�T�@��g-�s61�ݪ�ߛ��yU�P�����c��}ᬊ��o�?�^�%�����������z>�hK��K\�q�3-���o�=�U�+%���*�ỶuЃd�<YD��,}�K���Q�rRb28KT�Q����M��u�	��OS1V�$_��d$Ɖ+�Y�t�lpR�Z����
���]�~yUG�)a�/5�1OZy�ut�>��M��6V�NTz=��y3��m2�HPSL2����P����+$)X%��FFTB`%���x�m{����2 N	n� �ܯɦU������'\:�w؍L�ղ�9y�����;#s��@�]M�	��eI���H���{i�-��r�����FOU�R�t�I]��c�L9����I1�6�R���.�=a���dN77�;�q�S�.6�l_�gS%	D|�tg�+>�F�
(\0|6;u �;��\�Ry�dF� �����i�6�d�wm��wx��Fs�C� �{�⣸tj��ưE���T�`LMMR�-$�`� �W�����M)δ���g��z �?�ލ�	;���G�
S�`x�`�q��a��Ù�,Em@�9|I%כmI=(9�DH4߉E멸5���{E̻F�\�Kw.C:)\��dy����9�z��5'�=�y����uV�&nH<'�N��LS|$v@�����kހ͚�8�ڣ�<�����u%z4RᬢH�'�D\�`Z~f��m���4���+x6[bg̞��k�����bN�w�aM�u�}V�T�z�k�/��R�>���U�V�U�%t��^�S���OM���L�끊�@3�o*\Ƽ��������_�k��n�b�0�_����a��b�J���Ǧ�2��D����Ym�߈�G����z@�(������cNHɭ$ov��L֤��,��[s�ەNS�px�C�X#u�vU�U&5_}��C����pw-�u*��A�#��]��0c�A��0�m:_�� .US��g��"례��G�X�t�v��]A�_K�!�H���)Vp�a'a@�N��U	�r4���R΍mU(�lָ�@ȒJ���up��KO��$�)K�xf���=$�Ĩ	�W �}ȥ�؞S'$́��s��	����Vǡ�n�j�������^d�6�:���%oA(O�Sһ+w�ۆu0\gݧn�3/�.�׋����A>����a� Ŷ3��O�)Ѝx洫�Gֆ&��,��8D[���{�ل𳑺�x��j��QˀTK�@]CBV�<�?�<WE�<�u�o��f:փ��A?���w%����u�k;��vK���R�W-�l+`�#If؎!m=iM<�S�Ja!�hl���# dt\}���T��9��@y=fʇ����q
q9�@R� v��v�~���Sh�r�QΛ"��X���)����̞`6+"�.��<b�!����\��,�g���	L��I�ҝ�5���&~	y�����X���k~�#�v��_��������
Z����J��Vy��a�;�PI�y�4�<B�=�{���)5r,�"�����.�t�%�#��]��X���]�0(Ε��A���&��� �*����?�klT!wH�\M��wًע�3?�=�C�4���X.��\���>-��1\��R诬��~tC��4盚ɋ�#�P|A~
O��+�
��Dmvfڪ�w]	�nXH-���'��,�B1ħ��u���ӪMF[�|�8���`���ݥ�Ɩ�]= 6���8ۯR3��A��I"��x:dSަf�(����;�S�x�;����V�@5u�Xa�5K0]�^�Ў�Lg1��V����Z���@���<
�r�L۞^�D���L�c�`�
��馮_�{����2<��kd���[�����:����;�̖��F�k��i�?~׼�'�����l��%�Ζ�w�#B��CΌi�f�%�2t�:"+��YIh�/�3�y|�}Lar�Y�Z�1^�~�̘٥ֹ`�����0H,��F+'�R2W�oy����s-[�o�������)FS&������W��5���N`%DQ+ݧ�D |�&9Z^|����U���5qDx%�-�u?�������j���F�J�H�qJ�q9n�T�m�	r�-�$���z��F���ҁ�"�&_�{[ϯ9�Y�|Ã�fhj��b�w��5�6s��.? G�!�0'_N`�"��
Բ��Z�סE~���:�m��R:�Խ���3E!�e�������8�Rv��Dl7c�z�����$-�in�&�;� ��(�(���u�z`�)N��-�1Ef!�t��ɇ��@z7`���� y���> ��2��!�z�(G���1l���eT����Q�D���dV��״����B�����h���� 8�ts����Qkl۽�Q�X�YETN[]��M�]�N�k���LV�r� �m!�|��IJ���g����R9ѝ)�)����|���y "~oة/k-O,ۭ�L��gCq���m�	��#NS�C&%�>ŻC�����[�jj՜����*�b�&�z��uؚM�b�)��n��Q��f!eId�y�lH�����v��l�����rF$^�9/^>-��hGp���iCÚq�������h�Qv�[�|%����)����4/$D�x@��p~�d�[qE�C��Uc�'>�~~nZӺ�v�b��5|��J�
W~)X�r�H�U��1A�����[�5s��{�s]����mdmP~��|Fh�tT�ĺđ�O\�Hu�B����w=�P�� 	�X��w��@��g-��2�S���CKta�M��F�����)��k�-Vko�BA7^7]���Nj�P�(Q�)�"W9]E����4��!9�RD��%��vϧ��x���_��J���y�s�XI�	�y�F�s�Q���d!�D���DW�~�NJI�\�K���x���#R�30VYI�]���T!
6eVf�D�:3�+zF2�ݿ.׊45��zus��yӶB��
�?r+҇m�J]%UY����u/�����j��ŦtS�ǃA��n.}1L��ɝ�N��H*�~o�D-��_��nG���O_�ԇmt��Z;�8U��Utt�U�Įo��A 3mhd��8�;(m)к�N�=!��u��On�}\�zk���^�|�u���6R���`�eבG�F�x��^\
 �=�u}F-�id�Z`��]O�?,X9}�QmMw�\�fB�
���-X��p�}�5�*����c�l�2K�H	"e��݊Z��g[`�K�2 ���yN�5�	1_A^�a��&�{��S;{���G���t�h�)��|[^��`�K#QzqݿM�?g��đ��i�b/��@2 �����^��Z���]܅U�ظd�AZ4�Y�_3p-#���y�j���gO&�[k$��Θ6)�F�{��k�-YΉ)�6j�Ҙ���n��	X���eB��(GE(q�I�y�����8����Ea [MW)D�l��(��ه �A�w>$;�Ȑ�j~CCC�a}@­_��4�R��s.�>pÜ(�����0=�L�@ǄCޏw@O&[L����Ɲ��T��M����?jSb[�W���6P��c���$W�-fƝǥ�i���6{F���Q��?�n��+|������7L�OvEq��w�J�h�PuI�DD�o�6�T��:��
�R�Ìy���P���t,|��[^�<����d���?b��1�K����۽�?g�P*�N�YU�~�q<e�,*���l(����$3K$#4�%�~1Lf�YI����D���@{��R�5p�����\D�����{�5١���f2*�#RX1�ImՌ+C w2"�-,x���/����$�c#�*��Da��R={qy��iHe6#�v��nԱ��?-�rX��v�'R�GL��Ap�pmQ�F��N졑W�����LN�r!1��/ϩ�."�������ә���Oށ����V�X�O��n�%
$Fz(_��-��.����'�D����\���T��j�W��,?���a��U`@1���Wf���RI����;����L�gĎ�aD	-�RG�Ơ�`���4�f����:�Y_���gsQ��ߋ�dO���8�a֑��2N-���-��h�w1c�%)��F"�߶����<�T\��C��PK�;��M(�T��<�`ؚ(5����L�u� �/̇� ������5�3y��Ww�^L�^6Ճ�p�
�qk[�f��U��ͩ9^���)����w��!��3���ӞV�nҳ�cK��~�}��y��\/\�v���0F�Ǜ���cbjZk1˄�v 0���9�e�l.����Ѯ����bt��)��<�5�{:�r��������v%��"����]kZ�<}�i�ԌĿ|jGDc|����QE�g�Eа�hɯI>5 �^i�zG��JY���8詚^s�'VM�?^����z_��"�u�	 ���E2h<��N��i���g�Þ,Pѩ\��Ygn,�g�a��Gcw��l�p��b'Bi����7��k�����Z�c##t�i�_���7����^|���U-ܟܕ�������o?���	?N���{��(V�h�o���v��������HΊ+�]w���h��	����JY��UE(T��x�(��)$�{�T!j�߭�(��C��5F����c_�HӢ�♿wA��&�*_	��a�>#]��)~�J��ש�3����;����xUw��D�)Tx���⻶IG��sg:3M��jS99�[q�I?ܘ���E�?���${�^y��e�/�I��} SҒ2���Ɲ������_@���h�<���+!��BbF��	�������~g��m�TH����l"�6ɣ\Ǝ�4��r�����Ж����p
��ɯ�`	W87�]h�\�JY�zF����D�ăU$�S��5���)H���8�����G"���-:*�8�{'���=�d��U��_��<�h�I�]�)�^����VV��s���f�'�\�o�=���N��h��zk)�@�w��̻������a��/M�V�!U:��M�tOq��U��f{L��"��:���Y̨BY�18��E)�m�ש�&�I<���|���x#3��P	,��e���I9�����#�F`�?TD�Y����J(ӽ+]�l������\-2|0}��5=��#�˥�ҏ܉b\ٱ�{J�;/�S^�y��o���T�����?�a2����cI��H����b��C�R<G"7�N�i\��A�Op���̾~%Z���C�V_8�>����Y\^"9��l��gpH�,�gj�����懙l�{�)i\׈�'�	{�`W�����'[����cx�-}?ޖ��Tu\�l(H%@�H
ߦ픶L^��� _�DT��ʸ�@1�Oc�C�H%�5bG�@����fB 6���
�1��]�}��M�g���?�k�O��v@�M!�s���o �d�L�r����p>v�j.�F�}im6aK!"���oŘ���S�cF�H�"��a3�	�u��-1��V��"�)Y���_{C^��/D�{g���a'&sM�/eq}3��n�ywܮb��Q4q]��\2M��3�:oU��>ڞ�GV����`]vf��6,Y[���q4��$a�/��Ds")�^���[�� �b����u�{�D�}���&�۪3���S����(��=�/�P���fCB/>o�~���/��q���W�k��ԪF{TԸ*�a���ֹ]7�+p�nBQ�g\��
ZĊ�Y٪�f��V���N#�/^��p�<�5y���'���}��>+\�k�W����\������)v5?��pVK.Q$�f���A�T�n��Y�B$4lȚ��,�y"��fZn��i����h��7�����
����t��J��~�R�����p�펰�րS�b�t!�7����С���.�n�y�8��!��h�=��&.��W����)�5oH�XDg	�C�vY�n���X��X���jn�:2���o�E�����e7I�Ó%xt�b/�	4���-F���p1Y�>\EF�R�� �㣼u�ٍg��h�P̳a��8/]���_���Ѕ�����H��%Y1w�O�����GeB��,֓0q���.-Q����p�9a,%��P
�J����nU��!9����~&��,
�O.�ኹ39Aٕ�m�BE�Оr�c��U7��
Ҽ��o]����/�N���<����˩/�oEB:��p�Qv����?��<h��|ۊ�$��tY��J�|�jD�$��{.)޶��?�*�"�%I�fI8k�6�<���o&�Q��,
)�c�.�ػ*C���ꕸ`p����C��i߹��?���K����W��<������ޔ�(�ꐅ���0�|7����g��_|"���m�7go
����P���Գ��N�peC�O�L��Os�]e����9�hB�<��o�x��lRSC8E�	9n�r�罿y�:ť�"���z��Ƹ*^�)�.GFmY���/N)v�K�Mj@���L���Y@�ً�����w�Y��2�w����r�33Ih-y�� �DB���-�,)``���9�3,�V�s̭���
���,�1�4�	����D�ZQ�������믜�'C��>Be��`N����)����Y�k� �f��=�a��n�b7�NW�GL'[��mٻ��Ȣ�?�sgd؜�`�u>D}�� [ ��X��t���_ǳ\�JZ��d��NY�	�EbUCh�I�z������+xk����ű%G�+kc~�y�%v�3�\��G��A�Е�ƛ�#0 De�9X	���j2�;�ھ5����r��ZJ����-U�J�l�
��\���K�f��㐫چQLݐ=�co���>�;��,'j3������x�B"s����� 2��e��;�<��N�2ϗ��L3����Z�������J����x��$���~>���� ��C�7�u'�Z4~9�Ƈ�߆��FM�ָ�i�E�͟:J���W�{O���#�hң�W=F��/�փ�y)�D2����O�O��^d5�Ձ� Z�<���3S%�Wm�����DX�h�Pb�W1�!+��iN_HȦB��-J a���5[}C��\�嵱�<`��y���@�cFE��o����R~ܼ�.�j���=��
�@�5���1�g)�fl��s�c��NCH��q�Q�� Հ���}��&0I8h�����c�u�h��\i��ދ:|�u��I&dMc�<�"��8�P|��(<�+��s�;bg��,��4����YYh�]��A�^�%�B�2�����%�����j���_�G�����
5�BTo��vJ�IX�Lzkpo���S@��n5�����
��B�(I��������%`�x�"�|E��O���s�t<�����*�>�O��15�: E���e!T���.┬o��OS>�X���ͮe�?�"�(1���y+���X�}�n�qbG0+�Y�f�D�"��j��m�ލ<��bY��Z���SnT&���`��Tw pn�u���3�5/V�1r�]9�XrȮyN���I$�Pm,�˱��j��铔L�Q$����[J�q��@������U9��(S�%Sj(�������c�b~��S���3lL#N8E��1w��){�����-zy'�t�Z��߃�0u�z @,��<���(f-�	1�;����^�ݖz��u ��s�>v�3埚�Ԯ�	򭟉�����2�3y��Dc������T�$&n�~l�`V�e]�g7WX-�,��MR�!�
_�����^bH�ʃ2,�s�a�p$N�FP.�o |xb������������ ��-u
F�t��i�@�
���ô�7>/E)��ڷ�3:�Kv����bq����2^x��F�':I�������E]2$Ъ�kyx�ӝ������P^>�
�Sy"�|8C�����d��؅�GP<�EA���D��_����]D�`(�Jt�D�I�ҶQq��%���L1ChG2'���?nz5�1����ݽo%�Ea��i��!r8|EO�ڼ
��"�eD�b��2�0|1v�-� "<�RQu��k�-�0��hgiN��c�
�
-���/f���q����Y_ϓƄ� �h��r�I�8���EZhF�[PR��O���))>{ U�����;�z3����y�tq}�h��'�͚�A�� Iu;�l��cC4�������q�D��1ф��Ǒ;�7����X+���!!��fOx�8]����J�[%Z��pIb���>�j� ���DGV�yb������݃Y��7Z"���*@]5c�俁	���D�x�_xj+�F��=�ٌ������8vʾ��R���1B�޼b6�n/��c�Z}W��0�]�-®�	�#f�`�>�4M��Hǂ;i��A�B�4�lI���h6�9�}L�݌��c�f�ؠ������V jkD��u�#�[�Cw��"@�;�E�*�jD��B�G�nu-��=pװ�k���A�U�L]��DZ��g["�ۉϽ��99|�g+�Dc��]o�i� H`��Gu�>�F�����r����W� �V��ǹ�s��B�_���n�p�pԉ�e�Ey��m�E��X�z<�(?��>\ۂ�zET|H�Pk��1��5;XU���l�u�[�#�4^����/��곪�GNn�J"��|�/r�G�2�!_`�B5�a�D�Q�@�����,�۽���8���	9�u��&#�G�Y�&D�P�[>��m��m�t�~�g8Z�x	3�-�'�ױ�74��=G�>��`�H���1�!X!�/KH<��%��{OݑgE�;��m٫IMۡ�Y4E�[vO��-�1���.�,���=�9M���ߎ���gZ���vexzZ��/:��3Prh$��ɜ��'b����+�~����k0~u�ڃ�sL�0%�RH�����Kr��Vf-G��a�&5�D��gd���HB�A,��Æ�SFZ���L�+I;h{��r�!�>c�D�Y����s�$���L<��C���V2)�b�2��D$B��_os.�PR��]��0� ��G��_�c$A,h��;�f=c���8D��B浊�C�@�Yl�wt�Ek�60�B��G�c���u�y��'��Sw�^3Rc]�b{�U��"e?�����i,��k�I���$<�
g����g@9QJ�i���ό]n\jy=�2�R
���9�u?\�Sk�=4K���j�Ɨ�H��c�j�}��.�W�Q�y�?1O��p���e�~�@�,�Cy����ѯ���"�����:AO�՗�@No��[�,��u��-&۷��w5���ON����3%&&7[�q|Xd<r�s�hC^�=�>xD���4ɁX� ڏy��5X��wfs�򺑊�P�(���{����( �v����:��O������#~�o/��Z�a���_���c��Kn�����T�!��jxel�T��S��{"�C��~���?|�՞��.�W��c_�Ƒ�`hƲ��O@�0�!1���3=��@O2Y,�;�Fq/�KlF�e���a҆B�w�q:V��"V�]Gd%�$�D�A�W��&(}Y��QQf
?-L]-��i�R���a�� ��69�q%61Ų����gҿ�����s��9�XJ[w�ؚݹ雷pn�U\�'i#���>:K�P9g�`�
9���IO3�P���.���=�N>h�Ց0ży�ʄ/�=]?�f&o1W�ts�Sj���U(T��B�C�O�����G�;��x^0(�O�byu��5&L͞M\����q�a�[�5�Q����}T�^@�U���f�w��~�)yv�Cq$����J?�̵#���l�_���L����"�A�C�V1.��ZgeSU��-DhxQ�VGŇ��6��}ʭP+�{���_�A�أrl�:�4�����|M�p�,�>8���>E�w�pxs�7�������G=G�RB�+�
!�F��>?,�fU9���5������78zDX��r5K�N���a��`�4!���
+�i��O������������Ð[0ͺ�}��-�,�~�mq��x �[����%Qc&ݮa�����U��`v�~��[\�df6-�{���G
ܭ-��Ɂ��cl������.0�8�	���C�����[�#��k,HU����NT7��"l��#O���X)='�9u��)a5�Xv����ۓd����i��3	�I+:򠲹k�R������bY���[������ꌫ��[r=&�=��e����2�����SR5�h�5_
O�a�����o�b����-��>��MJ�_��!��g��*�(�f��n:N�GI'��v!9���R)�D�cFa��RNfD��7x�3�5�3��%60l�@�r��mz�%A��S+L(�� �՜�[������sA*���Q��v�.z��W`���ݍH>p�P��y�_4`0��M� T��LP ����������C���k�L`�`��֡��_n��,v�k
����(Ty��=��L�H����k����5�Y����Aኼ7���u��R��E���;FRk@m�tI��Ĳ��׵���t�'y ���/\2]��sT����_\T�P0��|_R+&^�G�$�ɼ�XU:FS~2?�d
?�i+4QY�Y�-���h�D���av���[V뫥�c�Cw]50�bzG�ơ�zK���w�@y�٠�6&�g�t�>��e�Mp$"�#�/�\�����JHL���V�G8|�pD��v�Te�ng�1�w(�F I!��:v���u:6�Z�"����H�`�/z#8i�	�B/��X	�,U��)ˠ�6kx�6uh�zU�t�h��gʭ~�q�zXDhʞ�J�C:�#����W�l��T+���?%?h	p���n.R����[ĥ\���la�;�n��1:\�f-O��+����d�T��:��0�4b^��8`9�������+D׈�v$1A����U���aU�g��NR���}ʄ9���d��bɅ��~�WsLsᯯ� pO��|�B��ء}[K���C�=�������lg���e �����rT�|��B��ů��j_})���t^)�����Ʈgq	$d���R<Z�w!p+�<Y��8]�w�ʖSG\)��7qH�.���&��H-R5�e#3�eO>�o�GM�:��Ӊ0j2b��yq9ӽC��q>{��d��®
�^C4Յ��4���+*;�Ue��H{�;z,��k��)�&��so�j-�oܥj̎�����}�HE9�89��9��\���єK� y|)'B�,�ˎϴ�C=@���=����s�B�WOtkR)�&t����p)���hV����+f�/K=�݋��&�V͞e�����ڣ��E�<٫����0[.�P�=bU7:C��q4�R&5�������obL'zPAAQ���d�ٶ7ɛ^�ݎ������7kN,5�22�r�P��V�T��cŧ�KQ"����Q��i�v�Q
5-��33=�oe�%~������U��ф����ڷ2<��=�_�\Q�QrA�����k!1�ޏ�o��[�d������GUoĨo�e���W�Uʏ�TV�w��h�ű������z��4Ykkܟ�]ZZ��M}m��{�)�
�ځ�Ͻc�MzZ�͙�y?rB|WJ\z��
���)ww�@��^`�J2͋f\������Ug$"��h{y�� E㠅���4Lv$�V����<�(�$\�y���)���?,�Z ��^8�?e��μG?��P��c|�ig`���ݫ�&��кLMVE�����&-I$|�Q�k�J�xp�v�]Į����`�����I���H"�ڿ9ᯁ!���k��������Xˁ2A��j4��y��;S#�B�S��2�!�x]}��<p�m5L�ﲼdH&�4w�������5kL�^��I{L
S$/��#��Q���[4d�84_��o�ъ��fi�qm�J�
���~�Z���Ǵ8Z�����%R�c��X�	x\���l�jp^�ǩ5��r�&OQ����U�����u֕��[�f�Fa�?�:�r֝�_��:/�ɑ[fH�o�@�]��;[�<oi5����!� J���9�M�
�h��OE��8mM�HI���|Pڶ>��*�mC�%]�L�;�ŕ��`a3�z�蘻t�m�B����}�n�P���߽Bd�n�I"�N�Oqv3Cp��i���fF�:jw<ё�.��q�khQ1z��w%�����e�tt8�O�"��62��$.�Ѻ�_�a�S^���{R���ނ#4h)�( �J�Z[��p~ċ!쌈����Ĭ���{a�w<��Acs���I�MHF3y3�S���(��
�"��+Jt��d:���!�e��|���I�N��
4��]_���qc�F��~\�?t0�d���tJ:��	��ZJ�7�FNQ��\���lT�V�S��-�'�mC���J,6�����a2�����bL��`%�K� 	8R5�@R�(��X-5Թ��:C�<�ѻ��텄��3�� ��pDAw1F�C�4D����KS��,ycL���i��'�y�	$n���~8��&(��4_Z#���ʩOHb�{J��DȖ��G�	��Ҧ�ߜW�h��ǤzJ���	
������V��G��R� s���\9J�kIêƤ��Z��[�r��a��B!�r���X�K���ػWBH��6��7d�G�<�l�y���<�め�Z�bҍ�,Y|��|�׼s��MZ���.�[Q�,� <�
/B=Bi���ݓ��H�e�<Q	8G����˻��-Բ?6��`��zSv�Jr�l_��!]���`�SLȯ�"��,w� :E��zR��<�ה�>ȳ| ���}).�)20�v�G��P��_Z5r�>z�y��;�j~s�r��|BL�m§�z$���Y����)���,�O�$�>#��¢�c�v�ck#�u>F��ONL[��t���"����eΆ���h��z�I�b��;-^^�Ё���d�t*��ऍ���t�2$.r�]M����%��u^�p݄Mi$��N����-^|n�^�2�aJ������zT�JR�[=uoF��%l�0t�*�F-��9 V���8a�cz��G��>[��h֠�?t��|���{��������Eی��]���|g��~������B���ʼ��������)Dz��ג�{@L�~�"ڵ4��$�.vŠ.l��y?*ĺ���[�|�Y���'˟���K`��SԷ��3�n��7��9��뭙z"�D�9���hr����Y��WA7W�Zq�3
/�}C�N�_��ʿ�*������2y�=p�4r�Qy�Ɵ
M��B�4�n�U5;떥�\�J�t_ÿ�Qn�pEt�'�`�U��K�����1it:���_�_.��˲,T�em���)?[����U(����a��Q�L��4̋l�'�z�U%C����>�W�7��qhȽէl�E��5������=N��eC6�q'U���aq����4�LA�N�ʴ�M�"S>�	��\�l�^�����t>0.�u�]?M5����D?;L�Y�2
Wm�,��Y�Լ�u���(QI�$dKV9���4S!BPWz�R�RTab�!�^4��<"�����.L>���X+�qKS�f���^����#�����ؗQ]����2F�M�-�@�I5wr�K�y�b�*��$g�B����Y(���Q#��:�L���誢e�l��E�Y�|�I�D��
�f��}H>셼K�i�V��ټ`�tH�*K�rb����"�y���]ƪ��V�Q��H!X��8�,����<߹��B�c4�#
�QYvߋ �F�\OQ^�Cu���#?%ސ��¢�HS�(~�9�6��b�߱��;���oa�q����r��wꌳ!��u���,/A�;b�x�w�H,���E(�pin�f�'�n�]�M2�Z����$������*L��D`3eM�CWjF�|ȼ��]��c�'>��H� E�5��e��u�7�-A}ԅ6W�M�]��Na��/��0}5�jBw 'A��D�O�w�OJc��ƔX���$���^yk.�z���nz����b��E�t����D�����y�{�T�6ɉ���lu/ ��p9։�u�Ю�G%օ�-�X��?G�`Q�,V���f���J�|k���m���}{K��6K�_/�#0f�'Ϟ����.�\��e����OrP�s���K�ڟj��(|N�7�"�M�I��FOpb*���`rE�=FX�3�ӡ	=���Q��Y'Չ� G6˧�E�ukE�VZ���KWj��;|$��7�8�]��W>�=byeo="><��M\�+ɡ�hx1׊�d��yea���m�J�_̸�r������ϟt�W��k^.iG7l/W���'R@�Wܥb�aeH��l�b��x�\��,Њ#_������u����Լ։�E�jG$)�]�,{(.�ݤ�N�},"�
�S������ ��L#10���ۃoOY����N�Q�\�*��U���C_F�c0:-z��S�i�8���x����#��%�l�mD�eo%�4GEc
&���kU�u���\��x!f�۶Z-��]�X��m]��}��R�2�!8�mhdB��$m�>����(ۯ��P��	�$����%H�x�7{MK�{���!�_8}�R����~�k	 � 9a@�(�E��3��"�`u/�mQa:�!ڧ����lh��L�e��+1:$BG�јA%J���dH�C@�S���'Yg�k}R�e�Df}W�ް����$:�~�+n~>\�/O&YI����{�K�K�򂼺��2g|;7��$�|���a�*<8��o�"���,���7��S)�Tޒzq��M�FX��̗ ��gm�XY�N�D���������S˶�"�U��K:�P��@�v�:���8؉��W�R��C/�Í��3���:�����
��n�,��:�1�'5��S��j 0Ex�-��j�;^l"J�]Bț��.k�o���i3�<�55f��-QcT8Me���j�,�'��]J��Q�[�t�	�q�Nj:�J��BO�#��w�N��i�d���=�qmF}U�Il�M5Ķ�h�O=��]�����M��>�Uh�3/63���os�|���J���M-�#*#S�{7v�}z��=|K�^���yXx;|�~�!L�U	�ON�:���g"B�����m���� �/��"*J�G[P�q�֩� ��1A��z��*sW��g�x۞Ð�.ܱY�[#(K@O�o�FsI?��d��<� 7�������\e֍0�[ ��\�>��L�l6q�1��VmQ͍Q��	�`j�]C���9����̙J��݈�fl��-��0����8��/%�~W��Y����A/q�E4� �꠩�v��t���?���m�	�;E�h�����mV����z��G��z͐Q����~��ʖ�b�.o"%�<?�!+�tE���Ny�|���fE�̇f[[��^~m=��h8�C���Uh�}�,J�a_%]UT����W�a@��Ȭ�;k��ϵ*�gO�5�?�'�7 3�l��O�ds��[{�	^�R�_p��=����)����F��&�^��^�������s7�6�Dh�FlOq��WJ�]ĩh�/����}�C+�S�7J�����>�Ph8�B�t]�kF��k;6R߄�g��������ӷ-\u���_��/����-+�i�C�F�ur���<~r� �J�m"�O��>D�ڡr��
lKXx���L��.ֲ���.������T���8HY%dZ_R}�&s�MqE��'	�7� vL/��L��U�3����}��<�/]+��}wʕ�D�<=�m�:�-���"5�E:(�?@;����S@��_#�ݓ��.]�;��a}���!+: �k���zo�ʨ�R�=ܖS�bw�b� Z���l,��w�+.���}B�nLi4�j����4�}�3��~PCe��JX�;�֒1�_��{��8�^�V�����	�ųD�3�	N���0�y�;�헞�=�|ݣ�;�/K���6yv��>}�P������%��[H�1�X�ak@]����/�ל:Vϋ�5�|�e�,Z-�3f�<Y�v�����ǖ�M"��gi��,����9�q,�H+V8��L"�����t�ξa�eb�������H�}SA�B!�&���Z���p{C0�Fdp��!`2F7�;�u�%�K�\^+��#U��E���I���Xr��C��Vl[W���'�r�Z�loݯ��;oR��eBb��OC�'�]p��L�}�貄M����_fv�KsZ_�,Ҿ#�m˝��[-���Qwǆ	9ƚ�+$n�W���@Q���o��À����9��6aPu͂�����5E���<1�{83�����)�>��I�n~�j �؝es�a�?\س���O�X�\uo�6�F�Ҵ��|�L��d�nc���Xs�姘-���B�Q�L�Vg���'��ҝ&�s������z}���17f:�Ȋ��8�u����$&�n�l�[�/��,?�.t7�g)�2�ZvD�v�l*�zC�%��0����p��	\�Ü3W�4:`K�ͼ�O�?�+iwD��H��/"�ȏ�������`���q)}��V`lb�5!g�
sE����e��O;�����zl���/æ� �`�T�G�fL�T��o&��>�\C�'��Y�gz�Yr+$ur4��q?lAN!��>o�&�Ws��"�6v$(3��%�p�x�^���Ͽ;�����^�H4���Y؁�<+fP7��w��>Y�O���1{�'���}�����D<l �{�	[��ΈFR0i� $�DK#�7[��M�;	X�4�Jb�R����%����}P�4K�h{���+*\"0csM����V�/��+���Yd��*����i�9�I硁�4�	ƥ�r�Ej)�y�����3!�A��մf�ë����^����RX@z9����ȵ)�ry+�u?)ɏ;�LP^{� A��w�z�HU<�;tc�^�b0�A��_ԇn�A`W��l=�)|�B�><���_�C�4tCw?;������<8���%'���2��	e��C��
���Kc� ��]���fy��B�Ϸ~ǝ}ΒЄh]<��Uo�&0���R���ْ�H^FRw�������>����l��8%��ue����P;~��j�-"Q��~�g<p�b�(F3�Pi3���WsQ������xK�VU4h�4�h�J�R�L�r��Fu� Ҽ����"깁�[��H��F����U%ҡc?�	��Ӗu�^2o�,�%�����x��d�;0��eج�H%ǚ2�GU����K�W�x�$<j�3JFi�p���:���^FLX�b�o)��0�~L{h�?th�$�4�U�.$�g���YB�o��TW��7�v�C�Q}�c��kZ��~��Dm'`�f2N=P��������?"=��z�/�~gQ����O�����H�-�
� @ p�Q�i�Q,�z}٫ޔBK-�+Yʠ	>��t���xW3B��'�3�
�ZQg)���6=�~|I4-7��_[j�d�Ae��{{���)ws���Xc���c�E�|��URJEu�a@���B������sT�C��K������J� U3-��MD��� a�,�+�؎!km�B���pxy�R{�p����������r��-�2�堅u�:���A}����]� V��u�G��%�|�Os��Vw����.���-b�~H�1�޼6��?�����ĭ�Wd҂�"����R�6��62��U������ӞKp�O���0��<���S������Pkl��W���c'k5�~Ü.��-�hj�lf/�&�f�lP0� ���ǣj�.dd�h�k����`����uM��H��&ޑE}��||�hx��3sN�=����h�����X3�A��Y:��Hǃ���C�z��pj�'�L|a�:�#t�Qt�ư�ġ����h�_w6�|�W�[�;�6���e?�g��Ɛ�c�(����w���F��tZ��I�>'�Y��a���R~��d�fWo�� �׵��Ml��5��G�V����a	�������H?�h����U�C	���߉3�&�6L?�M�٧���r��]!�k_����N�\��4{obP�9�'������.�$1���e2���D���$o� �)aȊ�
,f�������槁�%�\ȆO=��U�B�hq��c�(�/k��m���I��\��L��%��7���s���}�(�v��"N.)z$�L�Xx���V�.��8B��j����Q�U�>���~��~��B^��[��C�Ƨ~*��T�,3�xoZ�(�'�E\o���)#禍�b,T/��t_$�0a�'6�u<�jI@ҕ����^��ڡfƙ	&��^�����0x�G�;�2�Oo�M��D��f��R�ikd|��@8��D�5���.5AQ�8\�#��� ��/���$|����m�^"4 �7y�=�Ch�@�<�9��-
g]P�f L*�Dn0_ߓ�SE�m
x�WK(��&q~^��c(�P���H��!�.W��c�A�t�pD�ˉ����=-�̮ݟ��#QwVf�o��`���kah��j^o�6@�F��0�4��-
�f�����o~�y�T����2u<Lݥ����Z(!/�#"lWmk�[*���w�;� �uZE4o�� ���K�]1�g��B5�o����~���"SX�*sd�*Dی�4��Ď������J��v�k<-i�3���m�Ἵ���l��D����.i �b�Õ��+Z��^	~�C�1H��"���ۑ��~2��.K_ن�2�n���םOv��޳ݒ@S��v8�̔L��֭7G.vM��%T|���4_��h�����/.� u��IP��۷0{�S�@���-�֯(τ��j�wa�d�7��?}c��bNl�\�[F����k�� {�:������ʈ�1M�����Z���P�jVo�4��}UK/��1�D�#�+��ҷ �����
/ťw������w�12&>�F��(��L9������9��d�����'ںItv��ZTk�����bQ,�N��G�$�� �- �:R� �``*�f���C�4e�3�z�T�/s!��5�E6��=7W�B�b�P`��O��V"fa	Q��w`����R�u�?v�|?=b�ތI1^���8*�A��ť�k�M�h��#t)f����_����/�a���ڈ�|!����Q%�t��zs�����ez�I�p�x��FOEA⤠g�	 b��+�����ݥݒ��c���[Ֆ�����b��q���Z�#����e?�pL1`u��ֱ�s��$�J�c+d�� ��zR�����/�&�%�G��J�?��� ���H@�h�� <�G����M�o��*���8ͦ�T��]�U>�=MB�X0;$%��0uRA�=0�7ёW�U ���͝dK�nH�Ə����0������W�P���E���t���⤦�zy���$;�\kK��2��{��)A� ;^�l3иE�����y�ͣ��2��kp�nZ���q$bf���.ٲa,�A0=�۫�ӻ�����KaOȦ��Bx]cW������6��2܎�zJ�e'��7T�0���A[.���A�������R��j��]�KG� 	��+,�0�Zn��S'�H��V���?�rM#�\螱�&?�>0��V)s��$��\a~4+��,��h[��8�\[Ɔ�::Q�4p_��¹���踟�ٙ\K8�'-��K������7�D�I��š��ǿ�`g�ҺXE�0kF��+A�sO����u�T��kH���Ʊ��mv̗�k#)'l ��襺�&b��K]{&���3:3@>��8U?�Kq�GVG��U�fs��'��j��?����-�� �kO9���0�Һ�ޱ?�)p���T�4���t����߼Q>�*܎ک�X��'�<��
.�,�r᠈W3�A��H��;]t�;�����)�ƕ����P=d���u�m��Z��H�gXTۅB�v�Ǿ�X��E|���l�6� eE��}�C��:@ɡ�
�vUP�;#̩[�͗�
 R�_~�AG⹱��ߗS�PZS=d�!F�ႁm/�fɬX{W^��������B��� x�6�)I���W�-�I|�L+�?<�E�?40VҎ��S
��ҕ�rK��.�9u�Ű�גSm�5%a�<)b4ԡ	`�
#�n�����-�=��R��߆k�DA6�[�\\A�R��V��1a�)�TJǃC?�r��O�^{��A�D���O
�Gپ�{��(�ٺ�y��k���sB�5LdSsm/�7��/�~�#���/�3��U�H{��U�+��kʋ����& �o!&UuWvV��D���o�6-r�I�X�,�%��sM�9��\�t~*�~&1Z1E�j����4Q���!�JD��Ӹ1�)� ��4�V]3r4cR{��}��v'�b���f
؁y8�x�(���[�,* s�f�l�0����\RN�xr�Ե��"�&�)����{�ݖ��#�E1b={�}~�;|��6�`�~w\A��Y-�iZ)�#����~�ϫ4*L�V�?w`�@��Df�^-/�Ѓ�pȩ-*4#�gP5���vL�q�,u��)��Z����U�H)�S �&�RX��ԅ�D��ߎ�˗Z4� /!Ɨw��?f�| �>F�8�p�99)�������^�A��NW��Vy������q|�K:���
]��C1R2rn���`��0��2޵�C����=��z7����6�D^�ff`[j�G�
p�$�!�%�1�9�	�}�l?z���!��~+���H��-9fCۖ��8�����~���~~��� (���9|V&ó�c.��ki�2�6�����eyC�4AM���R��c���=K��Ұ�q�^�ib�_�jd{���7����C�'�y9iTH���FLO9;W;��Bd_	��"����#�������mr5�LԲ���;L`c��;I!��z.�D���:��G8��3�D���i����^54>��ZB椁r�
O�sF��m�.F2�["�ș����8�F "f�Kx��!����b�C�l��De�B��52�j\���Y7hמԔ�>�� �@�{�W�u|��ӓB.�^�0!����"�^�i��<w�v�|xzmf���m'l0߄�Fr�C����r���am<�[3ñ8�J���sM��@� P.������|��5R���"Q�Z�7�h�#~,1W����A��_�����9z^���[*�<�@x�@.YKr\o'!^�~��c��O���kf���n��^�%�� A�u�?�+w)u"����*>}��*�r���G�|r�w�8����5�Ǳi�4�� P�Ċ+�:�Ds��P���v�n������4�o�2����{��R�5������[�f�M���·'�"���G�e�
�*�\4�&\��/��|FY����(�=U2{�J$L���w!$�g���9�"��v���Y��TB��g=싕2@FD����|�DT"�U��2����D��k�}��YK�0�&[��3�7�,d����l��@]�+Lj_�%�Ĺ�Ƅ�����g	(����l8ɻM}�iG�(h!�z-G�V�+��L�x{9��x$M꛶��A�ɗI��3޸�C#��Q��֞v��Io�v�zJF>���l!������'�����}��
n�q��K�M�i��l�B	O�[/���-s���f?�q�%,>�qG�jDn�=̊CвI5��5^X�e�4�����>NbU�n㫞�s�3�J��X*^�l{^��^�������פ�!�Ʀ�"����)�Q��,�'QG�e��tY���hyLa�6���7�WU��?s�J���쑷és~�@\gQ�`2LxZ�M\�X�!��D�I8���|t5�{,x��{�)K<��'�v���n�	��sUs��5�i!z����#
�8�/�I=�7�7^�m��l(�;�`���Uf�@q���J/5�ֱ���:�7pöu�ʯ���63�d��3�~mrB&��m<�d�+߁A�TP�W.q�]}
����ĘEǩ �6z#��"����;=���.�{��4H����?����ܚ���T�;-[5���`<�韊���L������]�.A�9w(�GN��f�����"y�c��mMM3Je��a����~�ó|~��s⨬[��s�CNvG;+^6 Av'�#�x�)���p�W����I��c����_c�1���Q�B�x_M&>�O"�}w)�}�[JM^|�hm�br�`���@��J��f�I����$@��ԍRK �b�;� к�=-�u��q&^:s���q{ޥN�z��;�`g�)������bT��ڱ^Jk���&SC�Tcy�!�a^	�!�.�Vlộ�F�C�=�X�k�G���Y�<m3Ԏ��Wk��h�Q�h�IK�E�����~��;ƒC�\����4uV�V9���
���L߷EaDP�]Anש12�G���@�S�J,$�3��'S�0��ɢ\%.���D��Փ�[n/k��TF���_V��#.��;<��Ft��+w��H��Q�;!lL��^%5�e�"F0�n4(�K?fʻ2�'�ΪsY\���En������z�w�����b.4�ؚ�r��e9�yu�R���Ąrr�9a=L0�A�{��+^����g��,���pX1MFj�Li��(�f�T1w֧�Vz�����xU�yt;3�����24�ˡI��x�e�B�$�ގ���\-mB�?⿘�WY�Ҏ냺�z���ӈ�3�c���I�
.���톯_!S�@n;�q&�A����]������%�K;��H�zY���U�BG܂�0˃̃ik��Q�}Q���y��Q�J���d���V<���Jt^���,�+.���e�u�$��15��2;�r� tr���f,���B����Ln�t���\� O��h���"z��``�j���ܻ	ᤜ��W��/�?�@�_�����Cv����Bk>�q�1J�����U�T��$��P�k3�*���}1���b����O��V�&���"�v �~W��^���"ne�`�Ҿ[W��yM��U��\��@|��3�gAV�.����R�`�C΄V1�P/�����A��hg��~h�
�Y�L��y�eh2>���O�܏�hD�xxΒ�f�u�{sϢ��̿!�.Y��H����m ��@�p��� �4���c��mx��v�!�+)s�;e[ʹJA�̝���[2́���p��@����ik�'�x���b�"�j,uH�0�V�J^�ѼA�J�GJ��zd춻���ϐXz��*��jc�玂^�P?���v��e�)a��Q�J�s��D��zS�x
�#:�\�&�J���$�o��R���>Iø��v'Z�	*�\��2�ɼ0�������p��"�ʙ����L�c�Ş�6�����n'h��X^ل��I:1]�X��#h���w0w;�����8�0Rx���ѫF ������2�=��P��Bh�[����HnT���뻘�w�u��w#v�Qݤ�J��(R������B�߄;���/�,sKJN�L�������s�N������W)rQk��Ōb����/3	�HL(Z����kD�6՟H�U�>}C�4�V~�R���'��y$"*:<&���P��!�[`���ǅ�����Q�w6>a$/��@�|�6S[��G�&�Sd~�_Ӄ� ���!��Y�F&@���}ra�}��XR������RCX�f���(�eHkea��j"��N����?�����+��{���q�w糞��Hd[�L��(�WQ2�h��+�a._Z��_z�a3 >a �����`�l�Ih ��0���X��Bk|�����"���Ȏv�ȦE�_�A]��&��%�x��}�$r����%�m̱J{eQ[�}Uo� ��@�0=?!��M��'���*������L(��V�~KV1@�4�}�CEN���f���Q�����0�XA>��w���I'�fV��G|�2�lbĉ�o?��.i��@; h�,���N!c��. z8p�V����.�Nlb╺�4���z������|��H�5���0�M�8޸H4���W8��(y��Z�� xv<5�55*��d��G܎K<�Q`�S���`-�oǓj�Y1��z\�����@�~�����Ҳ@� ]W�i��8<�������|�fd�O>j6�CW��q!��RB������/QA��.�yq��
�b��3������$JÆ�~�S�V���o��Dw��\���`	dH6k�'hDۧ��(�}`b��k��[�X>fSn�" ꄰe�^f̉@����M�Q�Ԃ�ԥ�}h�)?��x���wˊ�	ͯt��L��q���췹?��$�фQ�<n���� $X�q���tE}5`����4J�*WS^7���-����}��;ޜ�|��CԈ��$��ׇ����n�{�J"�L��<ޥZN�B�ï��7uq��J�{�@+h�j2������~���5����}��pw�8:X�D���Rɀ��Z�������_�xgQ��4��#D��
���q}r%iA�)�5�y���,B"��46"8ȋh�R�%���]�F�XGٶ%(�_��-�$�웬����~�T	k�v�7�0/�B�#7�h���a"�q�*d�y��R�(i�;4(���u^�$�ﾏ���v�-Ε�`�^/o3J`&g�X}��5��RB�
*�M.��!��L)�$a��\I�oP�gpW7��Q�C SC�$�Ԛ*�u�\;h���T������] �{��m�A�߯�	o#dٕ�KarO\�]�� �tg�-@k�ܦhE؎�t�v�6����t��+��^��h�<�0��0"U�>��=u�k��eڎ�l���AAm�R:� �a����h���当����V:���B�7�[���n���f<�0>�9M�
����&�c��YO�V8�ѡ����3Ѓ(HR/$���kq�9���J1���Q�,��8�,9�Z}�K<�d�N�M�&��Ɠ�^�.�o�<Lۊ�3�����cC�e��
ō�����EG=��C�o�Nqp?r{��${���;�ბ ��J���O�is�?!�y`�q�z��y5M�X#(�VR	�??a�?�]m��J�7ihF��,�*4PAϰ_��o�SCz9�,,�"�X�N,U����)<"��b���~b�a�1
 �6�(;�6���Re�ŪE���	ꁞ]�S)ʁ"��e��|��Uq"3Ň��Fsz������ IF�,}�]�%�Pn�N��R�����+A�X��q�2��g�'B��h�����uj���̨v%n�v3��U�TS:���@O|�%��=ˣ����=��NGĩC�����.�:I�)�Q�+An�pj�@KaX���2/'�>yH2�B(B�ǳz��f6�$W*h7��<��؆��O�ť������mxjI-��I6}��CtlL�\�n��Y'�\����2.�^��-Uh%OM�2W[��M�̜��k	�,���r?�Z�4�|�R���]L���)��`MD`�1�qsJ|��K�B�66�A��5g| N`��6��ܢ�kS�/�cL�iB��[6>wc��W٫��/�$��JM��`\�j߬��?+����X�r�&���h��r�#<�f�O �)οKt�g��T1�E��d&� B���0g�K���	� Q�iG:�>b��կ���R�<:�
���	�?����2�p��?ۖ����5�_&֏x�*F�o�^���Ĕ�v-z�e�jH^�(��*�Z4�؈�t�G�s��^�D�A�k��\(����}�/�[/�״��>��an�8�e����<f�~���>P��~����R�B��@)�O�T������I�U�ܫEH�T��~�!����p.���ta�ICi��{��Z�O0�珯��&2J,_/��&rG��&$��D����w���N�P���[<Dj!��O��<�Ĩ7�[� W��E����m&����*���(\�<9���q� �vJ:P ���b�[��c�Jf�`%_ י���U���.����"z	�l�&�i�4X��la��e�g�������e+D)�q��m7�]�%�~<�a�I��UT��s!�o%���
�o�י�l�g��CPc�i�#�S�`϶3�4�B_�cpS������`��	��������:�e:>�カ@�H��=6т�>�Nu�~dɬ����a�M�vT��ر�!����F� !󋸉�_�����%�!��~�9R�)���ʹ�@5P[�+ۊ�Vu�q�G6w�-n�8{k���b%�x�茤H�$�)�{O�͜�����8"�{���֨����΂��Mrn�Eq��],�;���
�#�u�ϙ/ӏc���\����8�����p� �l�k�
��s
+�nK��0q:ښI|���j݄����;�^6���*�^}�ͅ������������K;4��v�l�hk�������(8}��Y<+��8lt�0zQg�*Mc���Ĥգ�\�/4�A�G>�0^�V�wY���r=66�V�x��ǼW��C�H��������]�X/�G��Ę��(��ܰ��7x9!�i6�е,8 �.ޅ�%S��S�O����4,Ո�#yu���SxWH�Ou�Uz�_#�qy��YԒ���p}����ǡR�M5�*�U���!Xϼs<M�Q�l9�V��Z�5����������y^U(mU��DʞŲ����G;j]F�^�¸E�16#b]s�>��4��ۭ���7/ƾ�+�Db��b+���2����dsH��.jӛ��
QK�To�1`�JHd����X[��i�uI�C�=�W���6�<c���w�	�ufY���0�o���1��W��kǥ�4��x'6L簽��/Q�an-h��T���8{}
�c��n�L�K��&ߠ�����������(��
��^���߳Z��W���ެ��/}�F�]���)8VD mp��&�7\���U &�Qnޮ��p����i`Ę��O��b�<�Ӄ�Y��C��r��g���*U�4_,D�u�S	�f�_��.c�69��}u�X>�ɀ��x�ee*�]:��	�;�EY�n|�k��qI� `Z��k�����(t"���Q[<���%zA���=S�����k��p�ՠmT�t����NBN��7.�h�K�Qum�S�R�
q�'E#�k�k�d�R�G�6�jDMI�Cf�cF�[�]�6+	� ��[YEm�~!���(Q^�-ݛ;O��hvr���W-K�ɜ���Ih%��}��L��ftr�ɹ�:8~�	]���
�''DT�����5pV-�{y�.KQۛRvW�j !E����ʦ�ϑ@��7��3��ꨈ�$�|�PtB^�y����k{�2~�mm��pfy10����7�.o��R ������n����=v���c��z@�f����bT
�:�DZ=�9Lh)�)!�Ȭ%[�
y�O�d~'[�6l�{4��1���N-ױ�0s+��i�o�xQJw��;�[�mF%��c��WO�u��_?@�=_����|�3G�Ǳ��Aݦ�y�m�j��j|�U���؞-tk�3�ܞ�:�ӡͦ׊��- �x���>L�{J���y�e�f�d��'��w����&��q���)��T���ܳ��df��L����%�G��E�U)}���:d�B�CO\Y��).<��L�5*�Q=�d��	�c�~(�z�V�ƣϙ,���>��+��鎁��"X��'���w��e$5�����1%�V���4�p��Sj�9��,�[4P5��٨����Sfzv!���\)�����\ V�$e≽m��z�
q3�91�I��#��f��*�Y���ML�Ȑug�O�����#�Ս��PZ���lL^DU��[N�ߞ���4��ֵ|+���;��JAweG�pr��+�-�z�dS�K�8�0t����G���a�<RYx�*
!� ����J�"y�j{u�F�i�	�}F�ƌ�ρC��X���g��y�w�N��R���<��zI�"�,��W�1LF�����o���v���� ��re&/vV]��Z�M�
�k��@�(z*��Q�	�s�@֍ǈU�HU�����\f������ױ�~]��Ӝ"N`�JޥB�ӣ��j��7�o�awZ�^�B#�H�+�hiB��
����J�5��08�'�mBI�2fY�<�D0
��uR�H%q~��fȞh
�#��q��jũ��^j �{� 5l?�����}��X�8��0��j��ա"��>��.�����0wa��PvC��6�M��PO�D�mt�b����d`��,����U�������������}�f-$���W�L�˒�TS"�q�P�����)�i�@s���#��K�x?_A��J��l�q�q�:FfVp,��*ր9 ��b���4j	p�8KΪz[����V�po�PFP)������Hٯ��nU͔O�$�+V��q�Cx���;�K��)ħ5P�f��M{��]����ߺ���!���B��A���)-�9�� �饟C���/��0���y�aA*^�~Oz$G=x�����,M���?����z���}Id)("��Ӑ�m?c������Ɉc����UE7$+.騟%M
�2>.��(���9{��l\?�,�����v;�X��f�/߷څ��Q�eO��!�U��g�E��v7��3V<Ǹ4�:˕� �]��m�ր�:��>:H#�4bUW�NÜ�:������}yBC?����>�Řˋw�?1w�Y�kȗ(Vqq����XI���e���)[���-��'@�(���J.��qV�s;Ae<����R+AZi�>@W�>�7��9H�fK�� ��
.���r���6eEKXl3�7a�Z���>�y�PW&�u[Q�VF,����E���+9�4�{��@"�V~�>ڊhd�xQ033��`�ˇ�IZ&���!��[�T�bc#�D
���K�u9nx(�%��tM5}� �GV /Wt}˾H}����h ����c��h���������)d��$��|8)m ���Al���9�q�t!�B�=��EC��(t��b�5[�[Q-�k��vr�˦<�)��[:X�.�4l�״��9"��P����z*��Nx�io��mǱ���-�J������|��AS0љƪT���b(N�?��e�+�vg@�ޘ�<|a)[UE6^�x1Ų��tigbft1�Na�"����Za�H��O��Gbb'[-@���Qf�3�?��� �9ڤ�H�BE�K��\^�u�2M�I0Y
�w'lǨ�n�Љ]^����a��XB�6�ⱘ��~ ���TM�g���y�:Tv�{�u �K��T�i�LzK����J����X� �BdX�GaߐT��9sit��g�+k�f��t�i����l�'�x ֜�~����gV�3�t�\_��9�8�Gi.���d�L�e���Pn׶�Ok:� �,��ݝ���iG\�4
�償(�am�Nyi�U&0��% -j0t�Oi
��]��uXɐq6E�;���܁<�B��LEb�Fo�G��ȼj���r�К��D�QrwZ?\�!�9|���9�{�/E=�ф|�-H��7ե�3�ݐ�(|LA3S@Z�CvK��Y��G�j?��2��� $g7�<+p1�SI���q(���p&Z�����b )B�g �u�
N=�:L@!{G�U��:C�k&�H#�P�v磛�S�]������K��ɍ,�1�k0���e/�3D�Aȗ��HƑ ��aE�7�f.��")�p�og��U��	��v3`��׃<Plq�~�]�
�`�$���qR9"�-H*]����]����g&tj���2�	��y&���̢U��/D�R�D^z����ʡ~ا�s��+�7��A6���,�Q�6� ��^��a|�l�T��4��T�Ty����v�S*�GF�Z��X[���I���@��I�v\Y�w�I��>q��*�\;k�5Ј\A5Ze���i���ν�Tc�}��/p��:ⰉE6��2�����P7&��1�͇w��B�_��j�����Õ@YC��Ӕ"��S�I���F������ұ�]���V�zZ�9-���|'��o�Ȑ�Y~�#��qS�^bq���5�c���(4�g�TL�,�,�-_���-��	7��y/��\���0&M[dJ��la���H��U�c�oO�i�KM̼�c�gf���*k���Y<Y#p@�3����vf巂��vr^tF
8,��S#t(�?�����r�k��4a�%���i��ћwӅ��!`���Ѥ�Ohz������f�
�j����Ԛ�RGݓ.d���	Yw��57�S��Ӫb)
�D�W�a\�~��3)�ҽ=��'���Z�<�Da�ݔ%�h��d�Lx莨M��H�ưr����&Z�<6@e�yVc�AԿy����_˳N^䠢�:�I�D�7/IR��4��۩rQ�e2,�ƞ_ˉ�F-�w�S�!�T�8�8�S�v�)��[�HdVVFpo"U��)�I&l�+ΰ�<��Q��� �{aG����Mt*F�S8��/�DO�ñj�Xu��a~��6~Ә|71 ���J*�~���Ve�����DAto"��E�� �]�mрv�ro"��l��q׎9��J	� 
b�)Y���:؎��B5��B�eau�X2�RX+U|zR^�F��lz"�(�>;,����wFK����!�d�[P�K�adP��}�ߥwz�#D'��� �S��/f���u�(��c�޿7�o���P762%�{^pZ�!]b]�t�0t�}!�
P>Ut ��f@��;�����u��l���y<|��H]9����n�1�^ղ�u��y���ʇB���,֌������̀���������"Ǫ>�KEg�Z�l�������,���bl�L����	d!&�]]�t+O�hw�c9�_��_�8�˱��.Z}�������ݵ�����+0�#��f#jl7�?�r(���RdX�鎰N:;�]�P����Ԕ3Y�p��;��٣S�<��`E�JK}������w���S�7���(P��ou:���V�s_�'p��u�׍��S �I�J�V����`LR��O��yp��ld�DN���������u�+��8��͸ff+&?�V����|�1&�ص�{��������K�G�ԝ��#�̸B�#{�8�Ws5���;��s��ڂ�&�}��+�r�˫�
���g��Ggζ������b?�x`�ِ�fLF�#���"�=�6��tqWj� e�g�����yJ;q� ~*Å�9����=)��㭝�����n�A���P��xE�:z�	*�����kZ˹H|s�"�b�����W�����f����P`����~ʩ�����EO�̽r��ƪ����B���P~����2W�Ε@�sL��#W�?��H4�ކ�u����T"�쏱ǀ�G�.�.�7�7�Gm �A� '���b��%��6�x��-��[;~��c���YBQ�"e�4�Y��j�w��B��p�������v�s��3��6~d�2S]z���=x�U#�}�w����,��L�Y�CQc��V����#g?lX[+J���XA+[r��BR#�N�(���d�7xK��:	0��zYتw���S�����%|:w �J�8R�
.�5����t��k�ߴi����5>�Yj	LtBd���K��c�_){�ĕ(���4wʴl���Z�G9U���?��X��Ψ����D��7o��8�A�_;Ō"I�f�gR�֥ :[GZh+0M�G��Z,j�VT]/hU��h��=��p-���G���[5��,(G~�2�y�#r���Aq����I,�
~z���4}XC��Ӣ���������l�ri��vXQ��H�w�� �*u)�p=T�ӿ�Hxb2��Q#�U��Vfyh��@�^
��i����-k��?��U��Z�s��.��2�G#$m�W�T��cT��2��Ta.~��V\�vҸh��i\h�Zc�ǫ�u���DW�Հ����>�^�Ȣ�z����Թ�ƣDgI��`Wg����T��K&���!~{|}�ڱ-���z��/�����=܀��ޙ�9J��d��t��s!)5U?&��6�yY�B�����~ߋS�y�Wu��췊n��)��:�}ɽM%�1�T��Z.��4���]ln]�6��kxxgU��iV" �0��$+��9#�,n2�i��=D���7�U�[���97����2__����ܵ��z��T����*��e��$�� cH]��yW��`��;&���@<��f.�N�#�[ �=�%� qkV�_���Ճhا7�����f2]S�����X�w�&�9��Vʟ����� �F�O�jӳr'��l4��y�Fvk�����jJS�ƈ-f��ta�;�"OE��U�2�~�l{ݯ��!�@�f"�x����䫫r�8aO�i=a1��t�=yy��~�:]R��R�)*�7��xک6���7U^��f!��T�Q a.~_ykB�&�������|Fl�3˼�n�;��<,����񢞵��P.�!������7/�D�Z�O'd���$N��H�_M���� ��.�blC,#�U�Α��v)*#[g\�ӣ'$�a8�Uzc/�;k	d�sߋ����,�4g�Z!Si��oo5�VѮ�+��dq�
��>na���������������6�|��Ե��p
����7�"^���-4��Ox.L�Ek
zKI	n,�ѐ­���L�l:�|xƆS�e��"G�8#�ޒ��]�^npP�������k��V�_w&��Fn�s�5J�/3��?��:���u����C��e�
d�|�oB)O��B6�P�F�!'���|ba.Hu�[e��@�E�hjZ9����I��
)9#���Q�e�u�B�%�E�;����>�,�oaH}�NG�8��DYGtPS�	H�t�2�X��� tp'
���!�M/�`����hݕ>���9�0B"
�]�i᱒$��(�YP��=eym�Z�7���.z�%�-n	�௝��L�p��,z� ����.�#�f��=N�.@�2�}��{�ِ� �k�[�6�@aJ�MT1N�י�YJ�BU���C��h�er��S/��UClw��o�r^��+!=�f�zh�.���"�_��Ja�W�c�|"��5{⩆�8�W�,F5KƂ��?�Lض����2Q#���|�����4հ��)y�>qY�*r�lOI#omP	�!rt�CH+~�df^
���Sy�����mp`,8h"R�T��L̠0TR�̽�e�s���GNA�e�{��ټQ��%>D}=�"Y��%�!�h)�i�{�r"	+�'����ڗ2�a��bW)�^C>~�U�j]���D�K�xK8�<rq�3�]�%�qDŻ�V���$�c �+� Z\��ҏ��ʣy�%ʃ��o]�h��H� �
���296��%�G_�$j�MɁ�Wf�NAQ,N
Vg�q�y�����s�K$C!B�C4�s[//��"ޗ:�*���3e4�����)zl�M���"��A�x��'�nIlC��:�^ǫ�����H{��"���xWC�d�N�3\����'��~��Fo�������������:�uj��9�a����W<��q���Tַ��n��0��0%�tǇ[�Mrn��x�h�Epԧǚ���a�B���H��"��Nf�g(������:�x���>���?�|�"��|P��F�GGR�4C�9*�C����DYdk:���'���|6�F؂�f}oi��\�ũ�� �(�T����7�i�kI�z>��,�[,E.=��ݫ��~�����C�Z�m@�
��0�	�H�q�6xh��DT�$��N�F��a�p�Ø��.m��	��G��\�3Ƚ"Ѭ:��}�1��L�]�@ΊH����|�o�ƭ�����d�mo*���B��j��W��}�rQS����Ǭ����z���S���FF�2e}1�|��&
U��3����.M��b�Q���Ԙz���@.�}�<8@���'�{^�+�W7�g�-RYOp��s+ȏ~��v�������r�y����[`}K�KK��2<��
Y�C9$���d�m��1��&t�O6$�+|k���iQ<PE��o�W� �����zbƽ�N��Q��lk�[J9������'uOUw�S� #�$�)��e� b�\�_�hT�@��������ă�TL��߼��C~^no:�v�>�/ 
�������!���6�{1�)Q@4�n����pu����}]ϯ�M�fC�x8KEf��Y]X����'����v������@���4���Ś�w��e���W�;k2{;b3.�`iPI���7I�%?�oK�d��>�|8,B�|M���3�|�Tƌ�$l�qM���b@(�gPY��X��ؕ�y���Y$�	�-
��oN`F���g�b@9XPcs�s�hq]J�G��>����H�.-m�.�O~�ʳ��i帳+��QH����b7�,�.Åj��[�,w���犵sK�k܄�HR���� �u��W��E�X?2?�h#�V/ψ;].����m�O/եT~Cګ��,�e�S�9H]v�8�	�}5��<��gE�(+��?&�×��{B�̙�M��.�w�i���Ul�4����Y��6-c�0ӷNΟ9+����v�#YA r)��u�3u��RxyJ��-P[�("�Q�3�-ݙj�3�H�+Fq2�o��E޴��u4�]�o�}�W���Hk*�XP��v�p���1�^5�������#�����f�f��sMu��Z��[4��y���%v1mjDi�v�W<����_��p�P���=?��J�k�ɏ�w�^��E�S��6�=�-�Nٖ+�I7x6ul6af B\?�%V�X�w/�<�CT١��1��B@u9Ϡr�q�����"4���m��%uC$�(2��A~��.ėy�����d��E"i8��a)�I���ҵ&�{�E�h{%�I�*O�HFf��� ���P�٠욆�+��wbx9��vQ~���!���\���׌\�	Nr^O2����~x���ш�Ty�ns�0�D��B���?��+�6�}}r*��Caa@ʧ:��WA�{�M8����(�G��iB�	�U#d�`S�����SěP&��-*j��LQY�3��Q_TG��Z��B�#kE���������������AY����R��9�:�\��'B�׌}�����ŗ>c��� T�^M�~g4��1���/����}׾����z�<�s��x��_]o��*��K^�^A���]h�i��?T���#�!�"�@�A�Á�c!��ص�"���ނ��Q`��{?�

�� �7�Ok54l=���:TZ�ڌ�.�笰j/@�<��y'e"*$C	�g�l��b�񅙨��q��yC�峚�d
�2T�خ��S8�ŴS@Y:C
\����kfs������f�)空�|n�@�T�E	�qи �jq�� ҹ���/�Y!Rt8���)VE��W��?���j��@)��죴���u�f�ED0������U�
�/�'b�3��/�t�r,��ן��s��oR�x��D	 �_m6Q�M~F�\񢹽ZO��-oć�4��^�gF�ޅfw5�:K��	Sv�C�l��Ch���V�>�Ω7�I_�0Ů"�TP��9�hoڞ��d�ȘxF��ȶ�� h�T/)�}��Ao�>�S�N���c��OYP����x`�Z�1�z�JiG�x�4�a��m��HV�ʏA�au#��J��?�1a6�:�M��;ܶΗ�X(�uȏ�e ��P_��3c�<ˑ}��V�4�Bг��1C,7����b@Ei�11wP~V��K̢ |��
�+�
{���Ǎ�.g���va]j���L�ȕ�9�oxE�[�zX�9v���.}��8s�M6� �����jeh[FFa�$��86�9��!���m	�2�/1d�ǖ"J �S����d��x�C��RQն7E��H{WZ3��S�y ����Œ���l^c0b����L��=��f=r��g��E3��:%i8���0�.#��v�f��;D
J��`c���#�̩d�"M$�8�IX���9c֒sۨ��Ag���U�یݤ�����������\�FG�����	i�BЉ�S>�A�U�<������8�8X�N"��xO�'�/���J 9�I��D	����h_�t�������$(+��ش�l�)b�
��G����	�˧>G���#��W�dX��!�P�˵[Sa��SZJ�u��(������K���@u�'�Gg���0��GP�e�YDQ�Ρ'���ѕ0��U���:Usw��������A=�4��K����#�bq�[p�*�*�z��./�2�'����;;�s^�_�t
�:f ��� }�Z�¹����N����w@�Ն�gŨ�����MDH�qa���zA8SQ���j(i=��x��F�C��Ԁ6����J�SAڍy&�^%s����_$mD$��d�����kF~~XԶ��ɟ.m1�|:�1Q��=T�[�(Á�0��{��J��YG��*��+��w���]�yiԛ��/	Z(�na�y��?���k���|��]���Wp�`7��D�v����z0n����λ�\�Ŗ��b�	�G�Kt@+�=���GtQS��(	��g��i�P�l���Ňt����5P���hϝ\&$-eeۘ�[E�<V$�=��B3�e�뷞j�pxO\�k�dWt���Lv.Jo�Y����N���~���i��%�.R���x��3�[��X��ꮠ�3h�3h���Y
�(�H�fY�^sM}:[<��tJJZ66���-��w�{�VC4?���u#���Ī�i)�c�X��#
V�璵H1vYt�~F���?�`ma3w4��SPMʩ�WL���z�0\S��Pb��rO�2��eD/ �iw.�C��ڥ1&{f��l.��i�`����������T�<�b��v`塴�RSy,M��C��H?�u��
��.K� �ؚ���1�H�G]S����z�KÔ6H��5� Ǥ��R��N���s�E�X����\�A:���
+�`�1��޶�L(~���2�I-��A>n�EYiT#�!W�����A� M@�8�?B��Ť�0{�젟������.�x8�a�}v�f��S>�P0��!��hP���ab ���d48��"a����qPX�?������L��15mW)^˭�iSo=5p}�2y����[�؜o��'���F���i1ED�S�@�02B�;AD�!��@vQ�A����:���OM"�=Y(1pO�ȲU����Z��
�����f�%1wxt3���=���hV��u��9�8T��c�wK*��o^�E���́
�p�5iG������wй�{ؗ�#�\��gb�l�;7e����r �]nw�&�~�WײE6�����o����f�r��S�rZ�c5�Ռ��묲5�']Gr��k&2ձ�WR!�/�%HLQjڌ_7�8����46sZ��'���	K���bs���q����%R"d�������_)C�����XMϛ WS��y�ϑ�����۹gO�x�B� 1�t8�"�C��P�P���<Kc�yQ�#�|CZ��T�pk�ծ����w3������㲈]������R�����2]|<��)9�"M.���1�/j��,��p��9�X�K߫���p�mIuo5M�d�ԣةI*ӭ6,����2�Ug��q�Y�U}�)�~1ܯR`�t���޹�,ȅ�>�=z�unr�@ba�x$��Hv��9�~cy��5j��n�R��8+��K|gZW"^�׌�e��=�ڦ�	��|�a0<)-&�^}�0�!_�]QX{�h,�������|��g������Ot�a�\CW�K7h5��?�R`\���g��_��	 ��th�B����A2�T��<i�E��1��,F�<e��.]�Z ��p1c|��Dı`���R}d��fF�3�ީ%���;3H�b��渕�^�v��¨97�N���{��9�4��(t�RƠ�m�%�*���%���=z���IML��^\-y�<�c���&���z�2�Lh`��Ko�;��Z#/U ���Ly,�翽���z/�X��J>�Ya�dZ�ҩ9��6}����z{UV�p�~����Q_~��aU;���?ꤎ��s�5��L�և��˾��3lɱ��] ��b��8[��2�e�V��A�ĝ)%0p�g��XV5#��Ė���<�,�5�v�����C�)��'0�l�����#�Hh\h��4��Ab�o�`���^[P�Bë�'r�^�3���A8��G�#'��N�0�2�ZVY�Woe�%��X{�s(0�w<���!9]����G�T����J��j�K����I0�M�AZQ�آ��G����5�g���K��Z�f��ޣx3
���hq�n�(������#�)���x�&�����̩��->
E3s��ʵ��x�S'ˠ����w<7�b�jp�@V�&Kl熺��N.41@<,���y���L@�	�A@������G��*܇�����~�b[��3Nj�$~�0
��w��oS�ǉ�޹�l�\[E��jn!D�@���A�����)b}�f���
�Y��W�[Hɺ�`�p|7�q���������bqQ��l��t�:�6!�c�7�?�#4ʔ��x�z�F1��x�I�b�/dHނ�l�������a�a�������8�і�ŧ�}�X���=�U�%�/���]9���u�=�|)�lM���,���w��Q,�r{U�������1��a��9v�j�a��.�E����'���H�ٱ@7���%�Xr�>�bX��N\���\�h�d���!"@�\���T=kUkX��*H�@�db���|D����t�^��zQ	q�lV��)���'��Y���V,0_g��4�$�����1�VU�X�ҼQ�V
�ᠠ4���.9��5kԾærP@�2��2�0q�T?���{OI�zR�-V�(����+��j�O�@�V\���y��[lwUyŔ�8�)I��7�2s\��"��vb�Y�鿚̭�ٽ2S�k87`�G�;Xqs����~�j%�)���a��߬&��Z�Kc��aN��z耕��Tx�w[�M��$B������]+8?(=V�z��eKT����Z.��G��Y���L�cq��k�>��!Ҍ�˫oW���%�3�U��#s�v��%���v�c�����q�N���J��/�Q���f�،Ӓ2�|/�",��=@
턣�11P����z�o�^!��hT���ą}ⶁ��Ƌ_n�UJFaSK?����*O�0q84���['���Ӓg>?h�Yj�<�
Yh:��4���p�����q�e�'��xջ�x��-;�H�ae�y�.T�*N�~m�;�� �Ɇ� 0'��K�\Lxގ._��|�����|���^��J�����0�}�+���\��!4�^���T��
OI.����"})뵸,J��HG*�C������_yM��O��g��r[7��m��&ui�&�"CSo[�����Q)��W�#��u��d���z�:؛r=At_h~�;þ]ͼ��N	8~r��Y�c�W�k���.*���g��#�n<�v�-��{|��B��.��ߌSy���������sU�kt��.�ɹ�\��W)ҫAnrfңT�� o��[�D��঄�E4D��z>�Kv䠢P��*ک����� �V�NE> �n�INn~o)(
����xNl�Zl>Nk�>ΰ��`�
~�x���:t(u5gp=|�(�S��T�ݦMgQqp���+��Y	�N�#��	龀,��)V��?c�F��[9`�/���-^���;�^�Ѭn=	ײ��b�9PP`+�w5�xfa�8����VG	�H�rm�����0�q�vp4MO'�OY�u*6-��4��H��W�K�*;@<zb�ua���G��nS�<?��K��f��k�By͔� �;T��z
��&'z� 6���(�@q�g�G}�-��F�}���d�	���P��4V�O��{�g���b�TR���k�-)3�����d���Af�/��x�US0���P~�O�컟0<�x��ț�[�)�0v�n=u��F��ȇC�߼-�G�G��|`�G`H�;K�;�A�ů
Ů�9�i��2��^��P�w��<I�A)�a�r�h+�!���'�����9�%O�pվ��_�s��
]g.�@��`1D���c�3{���^%��g�]���CY[)��)���<��flLA�3�{��!�F`l�lL��zy> v=]�]���w 2�>`g�b!B��QdE��h��UN+
K1<]�NKX!˨���p+�M0��C�>9��6�	����H5V�R�nZܾH��w�o@6�Z�@l�?���"�[������xK`�����`��}�k.Al��b������~G5<�x��?B�Zo4�c|�������NLzsE�`�֋37l���m`�l�2� ��8�$�� S)��g3���])L 
t$&�����˺䈸�UwTw�ml�m�j�&A�"�/Tƌ/��<�f�!�e�o1�=Edo�SHDJD�ԍj�9=��hN�\#.���k�Q~��2߉��	:�E�.�x6��C�U������Bo��(���G}��x	<� ���1�/�?jiag2���p�0#	I��Ǝ�G����ȴH�#��)1��UE�a��l�!��\7�Aب"&ۘ�����-5��VF��JY)a���R�U�s�ȕ�xJhe'=^�S��ӧ)��fƊC�=i�s:f� {��9�!���EO�c�"IzܺFw�����逗���	���hA�[�	��x��؜C�Y�E�,1��=:7lcN�U]�1מ<�U�;S�ȧ���8H� p���4���z���aW�E=�y��h��� A��<b�-�;Z��E������2��զ��mI������{��.����`�pp��T��ɶUYE]��T:���IoI�>�+�>2�"���)�wk?r�dQ4�K7ͫ;���誦���R�����@��(L=�L!�u[9P{�(���G=��t\'+����^�4�^S�ۤY��O��*��bz��'��	[S��wT��+���MTK���.�#H����/�7
�!�zM셬��4�j�R�M��˅�y4 ��@ϔ
���);�V�]�kuey���%�D��y!n�x�=%n? ?Y5���;�!���i��=������8S͉�Ҿ�Mj��CdSv���}�za ��\h�"�cs
Y�at��"HW�:����A�6�S1TO��ZSh�uZ��1��Yo���#���zZ&�7���_
0��H�_W��E{L[��P?ԗ�<��|kfD����0s}1��ݡ�g�C�.����{��ښqL��6�@��y-u@��֑�ſ�m@Tl5�y�R+�[�@�Q�B9}���]�j�(!C���x>�v���9T���݂ s|��ԭJ�h)$�L�i�_[�c����a�L�*;� �e��P��Jg7�7�I�/+�|Lh�K�����]�
�~�cՅ��,B��KPu�&�Ȟ(��mnܥ����z]B�o��2E�6��)���mK�H2�LAXUTJHpGf&���!$S��Ü#��.B��sh�p�;dG�8`����S�_��M�p:S�pV���/o�c�$QH/�~�婱'�>��d�VHՋ_�dz�K��%к>�v�Q���G��M��,\�o�ءS�܍�p?�s9t�
�"���[Xn'�{*���:��f���HkVg���J��ԝ��\�������R6�
R��MK���'>��vL��	�X�3��� 'ҝ�`����&���wԞ��,;j8B��ܔ�3�X\'
�u8Ԑ]�wZ�0t�%ֹ�y�"d^w.W����Ğ��Gd
11�넪�m�k�� *